5-I/P NAND GATE
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

.param width_P= {20*lambda}
.param width_N= {5*10*lambda}
    
Vdd	vdd	gnd	'SUPPLY'
va a gnd pulse 0 1.8 4ns 0ns 0ns 20ns 40ns
vb b gnd pulse 0 1.8 3ns 0ns 0ns 40ns 80ns
vc c gnd pulse 0 1.8 2ns 0ns 0ns 80ns 160ns
vd d gnd pulse 0 1.8 1ns 0ns 0ns 160ns 320ns
ve e gnd pulse 0 1.8 0ns 0ns 0ns 320ns 640ns
.option scale=0.09u


M1000 vo e a_56_n31# Gnd cmosn w=50 l=2
+  ad=250 pd=110 as=300 ps=112
M1001 vdd d vo vdd cmosp w=14 l=2
+  ad=238 pd=118 as=238 ps=118
M1002 a_56_n47# b a_56_n55# Gnd cmosn w=50 l=2
+  ad=300 pd=112 as=300 ps=112
M1003 vo a vdd vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_56_n31# d a_56_n39# Gnd cmosn w=50 l=2
+  ad=0 pd=0 as=300 ps=112
M1005 vo c vdd vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 a_56_n55# a gnd Gnd cmosn w=50 l=2
+  ad=0 pd=0 as=250 ps=110
M1007 a_56_n39# c a_56_n47# Gnd cmosn w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 vo e vdd vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 vdd b vo vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0

C0 vdd Gnd 2.25fF


.tran 0.1n 700n

.control
set hcopypscolor = 1
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=green
set color5=magenta
set color6=cyan
set color7=orange
run
plot v(a)+10 v(b)+8 v(c)+6 v(d)+4 v(e)+2 v(vo)
.endc

.end

