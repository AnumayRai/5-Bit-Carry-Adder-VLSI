magic
tech scmos
timestamp 1764415119
<< nwell >>
rect 6 40 163 101
rect 263 97 275 101
rect 230 57 326 97
rect 72 39 105 40
rect 230 20 254 57
rect 443 23 483 55
rect 4 -98 161 -37
rect 234 -97 274 -65
rect 332 -79 356 -42
rect 443 -74 483 -42
rect 70 -99 103 -98
rect 4 -239 161 -178
rect 263 -186 275 -182
rect 230 -226 326 -186
rect 70 -240 103 -239
rect 230 -263 254 -226
rect 440 -238 480 -206
rect 434 -312 474 -272
rect 4 -381 161 -320
rect 234 -380 274 -348
rect 335 -367 359 -330
rect 70 -382 103 -381
rect 434 -387 474 -347
rect 4 -568 161 -507
rect 263 -515 275 -511
rect 448 -512 488 -480
rect 230 -555 326 -515
rect 70 -569 103 -568
rect 230 -592 254 -555
rect 442 -586 482 -546
rect 4 -710 161 -649
rect 234 -709 274 -677
rect 335 -693 359 -656
rect 442 -676 482 -628
rect 70 -711 103 -710
rect 443 -766 483 -718
rect 450 -926 490 -894
rect 4 -1058 161 -997
rect 444 -1000 484 -960
rect 261 -1004 273 -1000
rect 228 -1044 324 -1004
rect 70 -1059 103 -1058
rect 228 -1081 252 -1044
rect 444 -1090 484 -1042
rect 2 -1199 159 -1138
rect 232 -1198 272 -1166
rect 334 -1178 358 -1141
rect 445 -1185 485 -1129
rect 68 -1200 101 -1199
rect 444 -1269 484 -1213
rect 449 -1421 489 -1389
rect 2 -1548 159 -1487
rect 260 -1494 272 -1490
rect 227 -1534 323 -1494
rect 443 -1495 483 -1455
rect 68 -1549 101 -1548
rect 227 -1571 251 -1534
rect 443 -1585 483 -1537
rect 2 -1689 159 -1628
rect 231 -1688 271 -1656
rect 334 -1664 358 -1627
rect 444 -1680 484 -1624
rect 68 -1690 101 -1689
rect 440 -1792 480 -1728
rect 437 -1885 477 -1821
rect 2 -2018 159 -1957
rect 68 -2019 101 -2018
<< ntransistor >>
rect 17 23 19 33
rect 47 23 49 33
rect 55 23 57 33
rect 110 19 112 29
rect 118 19 120 29
rect 150 22 152 32
rect 265 40 267 50
rect 288 34 290 44
rect 490 42 510 44
rect 490 34 510 36
rect 241 2 243 12
rect 490 -55 510 -53
rect 490 -63 510 -61
rect 281 -78 301 -76
rect 281 -86 301 -84
rect 15 -115 17 -105
rect 45 -115 47 -105
rect 53 -115 55 -105
rect 343 -97 345 -87
rect 108 -119 110 -109
rect 116 -119 118 -109
rect 148 -116 150 -106
rect 487 -219 507 -217
rect 487 -227 507 -225
rect 15 -256 17 -246
rect 45 -256 47 -246
rect 53 -256 55 -246
rect 108 -260 110 -250
rect 116 -260 118 -250
rect 148 -257 150 -247
rect 265 -243 267 -233
rect 288 -249 290 -239
rect 241 -281 243 -271
rect 481 -285 511 -283
rect 481 -293 511 -291
rect 481 -301 511 -299
rect 281 -361 301 -359
rect 481 -360 511 -358
rect 281 -369 301 -367
rect 481 -368 511 -366
rect 15 -398 17 -388
rect 45 -398 47 -388
rect 53 -398 55 -388
rect 346 -385 348 -375
rect 481 -376 511 -374
rect 108 -402 110 -392
rect 116 -402 118 -392
rect 148 -399 150 -389
rect 495 -493 515 -491
rect 495 -501 515 -499
rect 489 -559 519 -557
rect 15 -585 17 -575
rect 45 -585 47 -575
rect 53 -585 55 -575
rect 108 -589 110 -579
rect 116 -589 118 -579
rect 148 -586 150 -576
rect 265 -572 267 -562
rect 489 -567 519 -565
rect 288 -578 290 -568
rect 489 -575 519 -573
rect 241 -610 243 -600
rect 489 -641 529 -639
rect 489 -649 529 -647
rect 489 -657 529 -655
rect 489 -665 529 -663
rect 281 -690 301 -688
rect 281 -698 301 -696
rect 15 -727 17 -717
rect 45 -727 47 -717
rect 53 -727 55 -717
rect 346 -711 348 -701
rect 108 -731 110 -721
rect 116 -731 118 -721
rect 148 -728 150 -718
rect 490 -731 530 -729
rect 490 -739 530 -737
rect 490 -747 530 -745
rect 490 -755 530 -753
rect 497 -907 517 -905
rect 497 -915 517 -913
rect 491 -973 521 -971
rect 491 -981 521 -979
rect 491 -989 521 -987
rect 15 -1075 17 -1065
rect 45 -1075 47 -1065
rect 53 -1075 55 -1065
rect 108 -1079 110 -1069
rect 116 -1079 118 -1069
rect 148 -1076 150 -1066
rect 263 -1061 265 -1051
rect 491 -1055 531 -1053
rect 286 -1067 288 -1057
rect 491 -1063 531 -1061
rect 491 -1071 531 -1069
rect 491 -1079 531 -1077
rect 239 -1099 241 -1089
rect 492 -1142 542 -1140
rect 492 -1150 542 -1148
rect 492 -1158 542 -1156
rect 492 -1166 542 -1164
rect 279 -1179 299 -1177
rect 279 -1187 299 -1185
rect 492 -1174 542 -1172
rect 13 -1216 15 -1206
rect 43 -1216 45 -1206
rect 51 -1216 53 -1206
rect 345 -1196 347 -1186
rect 106 -1220 108 -1210
rect 114 -1220 116 -1210
rect 146 -1217 148 -1207
rect 491 -1226 541 -1224
rect 491 -1234 541 -1232
rect 491 -1242 541 -1240
rect 491 -1250 541 -1248
rect 491 -1258 541 -1256
rect 496 -1402 516 -1400
rect 496 -1410 516 -1408
rect 490 -1468 520 -1466
rect 490 -1476 520 -1474
rect 490 -1484 520 -1482
rect 13 -1565 15 -1555
rect 43 -1565 45 -1555
rect 51 -1565 53 -1555
rect 106 -1569 108 -1559
rect 114 -1569 116 -1559
rect 146 -1566 148 -1556
rect 262 -1551 264 -1541
rect 285 -1557 287 -1547
rect 490 -1550 530 -1548
rect 490 -1558 530 -1556
rect 490 -1566 530 -1564
rect 490 -1574 530 -1572
rect 238 -1589 240 -1579
rect 491 -1637 541 -1635
rect 491 -1645 541 -1643
rect 491 -1653 541 -1651
rect 278 -1669 298 -1667
rect 491 -1661 541 -1659
rect 491 -1669 541 -1667
rect 278 -1677 298 -1675
rect 345 -1682 347 -1672
rect 13 -1706 15 -1696
rect 43 -1706 45 -1696
rect 51 -1706 53 -1696
rect 106 -1710 108 -1700
rect 114 -1710 116 -1700
rect 146 -1707 148 -1697
rect 487 -1741 547 -1739
rect 487 -1749 547 -1747
rect 487 -1757 547 -1755
rect 487 -1765 547 -1763
rect 487 -1773 547 -1771
rect 487 -1781 547 -1779
rect 484 -1834 544 -1832
rect 484 -1842 544 -1840
rect 484 -1850 544 -1848
rect 484 -1858 544 -1856
rect 484 -1866 544 -1864
rect 484 -1874 544 -1872
rect 13 -2035 15 -2025
rect 43 -2035 45 -2025
rect 51 -2035 53 -2025
rect 106 -2039 108 -2029
rect 114 -2039 116 -2029
rect 146 -2036 148 -2026
<< ptransistor >>
rect 17 46 19 66
rect 25 46 27 66
rect 47 46 49 66
rect 55 46 57 66
rect 87 49 89 69
rect 110 62 112 82
rect 150 46 152 66
rect 265 63 267 83
rect 288 63 290 83
rect 241 26 243 46
rect 457 42 477 44
rect 457 34 477 36
rect 15 -92 17 -72
rect 23 -92 25 -72
rect 45 -92 47 -72
rect 53 -92 55 -72
rect 85 -89 87 -69
rect 108 -76 110 -56
rect 148 -92 150 -72
rect 343 -73 345 -53
rect 457 -55 477 -53
rect 457 -63 477 -61
rect 248 -78 268 -76
rect 248 -86 268 -84
rect 15 -233 17 -213
rect 23 -233 25 -213
rect 45 -233 47 -213
rect 53 -233 55 -213
rect 85 -230 87 -210
rect 108 -217 110 -197
rect 148 -233 150 -213
rect 265 -220 267 -200
rect 288 -220 290 -200
rect 454 -219 474 -217
rect 454 -227 474 -225
rect 241 -257 243 -237
rect 448 -285 468 -283
rect 448 -293 468 -291
rect 448 -301 468 -299
rect 15 -375 17 -355
rect 23 -375 25 -355
rect 45 -375 47 -355
rect 53 -375 55 -355
rect 85 -372 87 -352
rect 108 -359 110 -339
rect 148 -375 150 -355
rect 248 -361 268 -359
rect 346 -361 348 -341
rect 448 -360 468 -358
rect 248 -369 268 -367
rect 448 -368 468 -366
rect 448 -376 468 -374
rect 462 -493 482 -491
rect 462 -501 482 -499
rect 15 -562 17 -542
rect 23 -562 25 -542
rect 45 -562 47 -542
rect 53 -562 55 -542
rect 85 -559 87 -539
rect 108 -546 110 -526
rect 148 -562 150 -542
rect 265 -549 267 -529
rect 288 -549 290 -529
rect 456 -559 476 -557
rect 241 -586 243 -566
rect 456 -567 476 -565
rect 456 -575 476 -573
rect 456 -641 476 -639
rect 456 -649 476 -647
rect 456 -657 476 -655
rect 456 -665 476 -663
rect 15 -704 17 -684
rect 23 -704 25 -684
rect 45 -704 47 -684
rect 53 -704 55 -684
rect 85 -701 87 -681
rect 108 -688 110 -668
rect 148 -704 150 -684
rect 346 -687 348 -667
rect 248 -690 268 -688
rect 248 -698 268 -696
rect 457 -731 477 -729
rect 457 -739 477 -737
rect 457 -747 477 -745
rect 457 -755 477 -753
rect 464 -907 484 -905
rect 464 -915 484 -913
rect 458 -973 478 -971
rect 458 -981 478 -979
rect 458 -989 478 -987
rect 15 -1052 17 -1032
rect 23 -1052 25 -1032
rect 45 -1052 47 -1032
rect 53 -1052 55 -1032
rect 85 -1049 87 -1029
rect 108 -1036 110 -1016
rect 148 -1052 150 -1032
rect 263 -1038 265 -1018
rect 286 -1038 288 -1018
rect 239 -1075 241 -1055
rect 458 -1055 478 -1053
rect 458 -1063 478 -1061
rect 458 -1071 478 -1069
rect 458 -1079 478 -1077
rect 465 -1142 479 -1140
rect 465 -1150 479 -1148
rect 13 -1193 15 -1173
rect 21 -1193 23 -1173
rect 43 -1193 45 -1173
rect 51 -1193 53 -1173
rect 83 -1190 85 -1170
rect 106 -1177 108 -1157
rect 345 -1172 347 -1152
rect 465 -1158 479 -1156
rect 465 -1166 479 -1164
rect 146 -1193 148 -1173
rect 246 -1179 266 -1177
rect 246 -1187 266 -1185
rect 465 -1174 479 -1172
rect 464 -1226 478 -1224
rect 464 -1234 478 -1232
rect 464 -1242 478 -1240
rect 464 -1250 478 -1248
rect 464 -1258 478 -1256
rect 463 -1402 483 -1400
rect 463 -1410 483 -1408
rect 457 -1468 477 -1466
rect 457 -1476 477 -1474
rect 457 -1484 477 -1482
rect 13 -1542 15 -1522
rect 21 -1542 23 -1522
rect 43 -1542 45 -1522
rect 51 -1542 53 -1522
rect 83 -1539 85 -1519
rect 106 -1526 108 -1506
rect 146 -1542 148 -1522
rect 262 -1528 264 -1508
rect 285 -1528 287 -1508
rect 238 -1565 240 -1545
rect 457 -1550 477 -1548
rect 457 -1558 477 -1556
rect 457 -1566 477 -1564
rect 457 -1574 477 -1572
rect 464 -1637 478 -1635
rect 13 -1683 15 -1663
rect 21 -1683 23 -1663
rect 43 -1683 45 -1663
rect 51 -1683 53 -1663
rect 83 -1680 85 -1660
rect 106 -1667 108 -1647
rect 345 -1658 347 -1638
rect 464 -1645 478 -1643
rect 464 -1653 478 -1651
rect 146 -1683 148 -1663
rect 245 -1669 265 -1667
rect 464 -1661 478 -1659
rect 464 -1669 478 -1667
rect 245 -1677 265 -1675
rect 454 -1741 474 -1739
rect 454 -1749 474 -1747
rect 454 -1757 474 -1755
rect 454 -1765 474 -1763
rect 454 -1773 474 -1771
rect 454 -1781 474 -1779
rect 451 -1834 471 -1832
rect 451 -1842 471 -1840
rect 451 -1850 471 -1848
rect 451 -1858 471 -1856
rect 451 -1866 471 -1864
rect 451 -1874 471 -1872
rect 13 -2012 15 -1992
rect 21 -2012 23 -1992
rect 43 -2012 45 -1992
rect 51 -2012 53 -1992
rect 83 -2009 85 -1989
rect 106 -1996 108 -1976
rect 146 -2012 148 -1992
<< ndiffusion >>
rect 16 23 17 33
rect 19 23 20 33
rect 46 23 47 33
rect 49 23 50 33
rect 54 23 55 33
rect 57 23 58 33
rect 109 19 110 29
rect 112 19 113 29
rect 117 19 118 29
rect 120 19 121 29
rect 149 22 150 32
rect 152 22 153 32
rect 264 40 265 50
rect 267 40 268 50
rect 287 34 288 44
rect 290 34 291 44
rect 490 44 510 45
rect 490 41 510 42
rect 490 36 510 37
rect 490 33 510 34
rect 240 2 241 12
rect 243 2 244 12
rect 490 -53 510 -52
rect 490 -56 510 -55
rect 490 -61 510 -60
rect 490 -64 510 -63
rect 281 -76 301 -75
rect 281 -79 301 -78
rect 281 -84 301 -83
rect 281 -87 301 -86
rect 14 -115 15 -105
rect 17 -115 18 -105
rect 44 -115 45 -105
rect 47 -115 48 -105
rect 52 -115 53 -105
rect 55 -115 56 -105
rect 342 -97 343 -87
rect 345 -97 346 -87
rect 107 -119 108 -109
rect 110 -119 111 -109
rect 115 -119 116 -109
rect 118 -119 119 -109
rect 147 -116 148 -106
rect 150 -116 151 -106
rect 487 -217 507 -216
rect 487 -220 507 -219
rect 487 -225 507 -224
rect 487 -228 507 -227
rect 14 -256 15 -246
rect 17 -256 18 -246
rect 44 -256 45 -246
rect 47 -256 48 -246
rect 52 -256 53 -246
rect 55 -256 56 -246
rect 107 -260 108 -250
rect 110 -260 111 -250
rect 115 -260 116 -250
rect 118 -260 119 -250
rect 147 -257 148 -247
rect 150 -257 151 -247
rect 264 -243 265 -233
rect 267 -243 268 -233
rect 287 -249 288 -239
rect 290 -249 291 -239
rect 240 -281 241 -271
rect 243 -281 244 -271
rect 481 -283 511 -282
rect 481 -286 511 -285
rect 481 -291 511 -290
rect 481 -294 511 -293
rect 481 -299 511 -298
rect 481 -302 511 -301
rect 281 -359 301 -358
rect 481 -358 511 -357
rect 281 -362 301 -361
rect 281 -367 301 -366
rect 281 -370 301 -369
rect 481 -361 511 -360
rect 481 -366 511 -365
rect 14 -398 15 -388
rect 17 -398 18 -388
rect 44 -398 45 -388
rect 47 -398 48 -388
rect 52 -398 53 -388
rect 55 -398 56 -388
rect 345 -385 346 -375
rect 348 -385 349 -375
rect 481 -369 511 -368
rect 481 -374 511 -373
rect 481 -377 511 -376
rect 107 -402 108 -392
rect 110 -402 111 -392
rect 115 -402 116 -392
rect 118 -402 119 -392
rect 147 -399 148 -389
rect 150 -399 151 -389
rect 495 -491 515 -490
rect 495 -494 515 -493
rect 495 -499 515 -498
rect 495 -502 515 -501
rect 489 -557 519 -556
rect 14 -585 15 -575
rect 17 -585 18 -575
rect 44 -585 45 -575
rect 47 -585 48 -575
rect 52 -585 53 -575
rect 55 -585 56 -575
rect 107 -589 108 -579
rect 110 -589 111 -579
rect 115 -589 116 -579
rect 118 -589 119 -579
rect 147 -586 148 -576
rect 150 -586 151 -576
rect 264 -572 265 -562
rect 267 -572 268 -562
rect 489 -560 519 -559
rect 489 -565 519 -564
rect 287 -578 288 -568
rect 290 -578 291 -568
rect 489 -568 519 -567
rect 489 -573 519 -572
rect 489 -576 519 -575
rect 240 -610 241 -600
rect 243 -610 244 -600
rect 489 -639 529 -638
rect 489 -642 529 -641
rect 489 -647 529 -646
rect 489 -650 529 -649
rect 489 -655 529 -654
rect 489 -658 529 -657
rect 489 -663 529 -662
rect 489 -666 529 -665
rect 281 -688 301 -687
rect 281 -691 301 -690
rect 281 -696 301 -695
rect 281 -699 301 -698
rect 14 -727 15 -717
rect 17 -727 18 -717
rect 44 -727 45 -717
rect 47 -727 48 -717
rect 52 -727 53 -717
rect 55 -727 56 -717
rect 345 -711 346 -701
rect 348 -711 349 -701
rect 107 -731 108 -721
rect 110 -731 111 -721
rect 115 -731 116 -721
rect 118 -731 119 -721
rect 147 -728 148 -718
rect 150 -728 151 -718
rect 490 -729 530 -728
rect 490 -732 530 -731
rect 490 -737 530 -736
rect 490 -740 530 -739
rect 490 -745 530 -744
rect 490 -748 530 -747
rect 490 -753 530 -752
rect 490 -756 530 -755
rect 497 -905 517 -904
rect 497 -908 517 -907
rect 497 -913 517 -912
rect 497 -916 517 -915
rect 491 -971 521 -970
rect 491 -974 521 -973
rect 491 -979 521 -978
rect 491 -982 521 -981
rect 491 -987 521 -986
rect 491 -990 521 -989
rect 14 -1075 15 -1065
rect 17 -1075 18 -1065
rect 44 -1075 45 -1065
rect 47 -1075 48 -1065
rect 52 -1075 53 -1065
rect 55 -1075 56 -1065
rect 107 -1079 108 -1069
rect 110 -1079 111 -1069
rect 115 -1079 116 -1069
rect 118 -1079 119 -1069
rect 147 -1076 148 -1066
rect 150 -1076 151 -1066
rect 262 -1061 263 -1051
rect 265 -1061 266 -1051
rect 491 -1053 531 -1052
rect 285 -1067 286 -1057
rect 288 -1067 289 -1057
rect 491 -1056 531 -1055
rect 491 -1061 531 -1060
rect 491 -1064 531 -1063
rect 491 -1069 531 -1068
rect 491 -1072 531 -1071
rect 491 -1077 531 -1076
rect 491 -1080 531 -1079
rect 238 -1099 239 -1089
rect 241 -1099 242 -1089
rect 492 -1140 542 -1139
rect 492 -1143 542 -1142
rect 492 -1148 542 -1147
rect 492 -1151 542 -1150
rect 492 -1156 542 -1155
rect 492 -1159 542 -1158
rect 492 -1164 542 -1163
rect 279 -1177 299 -1176
rect 279 -1180 299 -1179
rect 279 -1185 299 -1184
rect 492 -1167 542 -1166
rect 492 -1172 542 -1171
rect 492 -1175 542 -1174
rect 279 -1188 299 -1187
rect 12 -1216 13 -1206
rect 15 -1216 16 -1206
rect 42 -1216 43 -1206
rect 45 -1216 46 -1206
rect 50 -1216 51 -1206
rect 53 -1216 54 -1206
rect 344 -1196 345 -1186
rect 347 -1196 348 -1186
rect 105 -1220 106 -1210
rect 108 -1220 109 -1210
rect 113 -1220 114 -1210
rect 116 -1220 117 -1210
rect 145 -1217 146 -1207
rect 148 -1217 149 -1207
rect 491 -1224 541 -1223
rect 491 -1227 541 -1226
rect 491 -1232 541 -1231
rect 491 -1235 541 -1234
rect 491 -1240 541 -1239
rect 491 -1243 541 -1242
rect 491 -1248 541 -1247
rect 491 -1251 541 -1250
rect 491 -1256 541 -1255
rect 491 -1259 541 -1258
rect 496 -1400 516 -1399
rect 496 -1403 516 -1402
rect 496 -1408 516 -1407
rect 496 -1411 516 -1410
rect 490 -1466 520 -1465
rect 490 -1469 520 -1468
rect 490 -1474 520 -1473
rect 490 -1477 520 -1476
rect 490 -1482 520 -1481
rect 490 -1485 520 -1484
rect 12 -1565 13 -1555
rect 15 -1565 16 -1555
rect 42 -1565 43 -1555
rect 45 -1565 46 -1555
rect 50 -1565 51 -1555
rect 53 -1565 54 -1555
rect 105 -1569 106 -1559
rect 108 -1569 109 -1559
rect 113 -1569 114 -1559
rect 116 -1569 117 -1559
rect 145 -1566 146 -1556
rect 148 -1566 149 -1556
rect 261 -1551 262 -1541
rect 264 -1551 265 -1541
rect 284 -1557 285 -1547
rect 287 -1557 288 -1547
rect 490 -1548 530 -1547
rect 490 -1551 530 -1550
rect 490 -1556 530 -1555
rect 490 -1559 530 -1558
rect 490 -1564 530 -1563
rect 490 -1567 530 -1566
rect 490 -1572 530 -1571
rect 490 -1575 530 -1574
rect 237 -1589 238 -1579
rect 240 -1589 241 -1579
rect 491 -1635 541 -1634
rect 491 -1638 541 -1637
rect 491 -1643 541 -1642
rect 491 -1646 541 -1645
rect 491 -1651 541 -1650
rect 278 -1667 298 -1666
rect 278 -1670 298 -1669
rect 491 -1654 541 -1653
rect 491 -1659 541 -1658
rect 491 -1662 541 -1661
rect 491 -1667 541 -1666
rect 278 -1675 298 -1674
rect 278 -1678 298 -1677
rect 344 -1682 345 -1672
rect 347 -1682 348 -1672
rect 491 -1670 541 -1669
rect 12 -1706 13 -1696
rect 15 -1706 16 -1696
rect 42 -1706 43 -1696
rect 45 -1706 46 -1696
rect 50 -1706 51 -1696
rect 53 -1706 54 -1696
rect 105 -1710 106 -1700
rect 108 -1710 109 -1700
rect 113 -1710 114 -1700
rect 116 -1710 117 -1700
rect 145 -1707 146 -1697
rect 148 -1707 149 -1697
rect 487 -1739 547 -1738
rect 487 -1742 547 -1741
rect 487 -1747 547 -1746
rect 487 -1750 547 -1749
rect 487 -1755 547 -1754
rect 487 -1758 547 -1757
rect 487 -1763 547 -1762
rect 487 -1766 547 -1765
rect 487 -1771 547 -1770
rect 487 -1774 547 -1773
rect 487 -1779 547 -1778
rect 487 -1782 547 -1781
rect 484 -1832 544 -1831
rect 484 -1835 544 -1834
rect 484 -1840 544 -1839
rect 484 -1843 544 -1842
rect 484 -1848 544 -1847
rect 484 -1851 544 -1850
rect 484 -1856 544 -1855
rect 484 -1859 544 -1858
rect 484 -1864 544 -1863
rect 484 -1867 544 -1866
rect 484 -1872 544 -1871
rect 484 -1875 544 -1874
rect 12 -2035 13 -2025
rect 15 -2035 16 -2025
rect 42 -2035 43 -2025
rect 45 -2035 46 -2025
rect 50 -2035 51 -2025
rect 53 -2035 54 -2025
rect 105 -2039 106 -2029
rect 108 -2039 109 -2029
rect 113 -2039 114 -2029
rect 116 -2039 117 -2029
rect 145 -2036 146 -2026
rect 148 -2036 149 -2026
<< pdiffusion >>
rect 16 46 17 66
rect 19 46 20 66
rect 24 46 25 66
rect 27 46 28 66
rect 46 46 47 66
rect 49 46 50 66
rect 54 46 55 66
rect 57 46 58 66
rect 86 49 87 69
rect 89 49 90 69
rect 109 62 110 82
rect 112 62 113 82
rect 149 46 150 66
rect 152 46 153 66
rect 264 63 265 83
rect 267 63 268 83
rect 287 63 288 83
rect 290 63 291 83
rect 240 26 241 46
rect 243 26 244 46
rect 457 44 477 45
rect 457 41 477 42
rect 457 36 477 37
rect 457 33 477 34
rect 14 -92 15 -72
rect 17 -92 18 -72
rect 22 -92 23 -72
rect 25 -92 26 -72
rect 44 -92 45 -72
rect 47 -92 48 -72
rect 52 -92 53 -72
rect 55 -92 56 -72
rect 84 -89 85 -69
rect 87 -89 88 -69
rect 107 -76 108 -56
rect 110 -76 111 -56
rect 147 -92 148 -72
rect 150 -92 151 -72
rect 248 -76 268 -75
rect 342 -73 343 -53
rect 345 -73 346 -53
rect 457 -53 477 -52
rect 457 -56 477 -55
rect 457 -61 477 -60
rect 457 -64 477 -63
rect 248 -79 268 -78
rect 248 -84 268 -83
rect 248 -87 268 -86
rect 14 -233 15 -213
rect 17 -233 18 -213
rect 22 -233 23 -213
rect 25 -233 26 -213
rect 44 -233 45 -213
rect 47 -233 48 -213
rect 52 -233 53 -213
rect 55 -233 56 -213
rect 84 -230 85 -210
rect 87 -230 88 -210
rect 107 -217 108 -197
rect 110 -217 111 -197
rect 147 -233 148 -213
rect 150 -233 151 -213
rect 264 -220 265 -200
rect 267 -220 268 -200
rect 287 -220 288 -200
rect 290 -220 291 -200
rect 454 -217 474 -216
rect 454 -220 474 -219
rect 454 -225 474 -224
rect 454 -228 474 -227
rect 240 -257 241 -237
rect 243 -257 244 -237
rect 448 -283 468 -282
rect 448 -286 468 -285
rect 448 -291 468 -290
rect 448 -294 468 -293
rect 448 -299 468 -298
rect 448 -302 468 -301
rect 14 -375 15 -355
rect 17 -375 18 -355
rect 22 -375 23 -355
rect 25 -375 26 -355
rect 44 -375 45 -355
rect 47 -375 48 -355
rect 52 -375 53 -355
rect 55 -375 56 -355
rect 84 -372 85 -352
rect 87 -372 88 -352
rect 107 -359 108 -339
rect 110 -359 111 -339
rect 147 -375 148 -355
rect 150 -375 151 -355
rect 248 -359 268 -358
rect 345 -361 346 -341
rect 348 -361 349 -341
rect 448 -358 468 -357
rect 448 -361 468 -360
rect 248 -362 268 -361
rect 248 -367 268 -366
rect 248 -370 268 -369
rect 448 -366 468 -365
rect 448 -369 468 -368
rect 448 -374 468 -373
rect 448 -377 468 -376
rect 462 -491 482 -490
rect 462 -494 482 -493
rect 462 -499 482 -498
rect 462 -502 482 -501
rect 14 -562 15 -542
rect 17 -562 18 -542
rect 22 -562 23 -542
rect 25 -562 26 -542
rect 44 -562 45 -542
rect 47 -562 48 -542
rect 52 -562 53 -542
rect 55 -562 56 -542
rect 84 -559 85 -539
rect 87 -559 88 -539
rect 107 -546 108 -526
rect 110 -546 111 -526
rect 147 -562 148 -542
rect 150 -562 151 -542
rect 264 -549 265 -529
rect 267 -549 268 -529
rect 287 -549 288 -529
rect 290 -549 291 -529
rect 456 -557 476 -556
rect 456 -560 476 -559
rect 240 -586 241 -566
rect 243 -586 244 -566
rect 456 -565 476 -564
rect 456 -568 476 -567
rect 456 -573 476 -572
rect 456 -576 476 -575
rect 456 -639 476 -638
rect 456 -642 476 -641
rect 456 -647 476 -646
rect 456 -650 476 -649
rect 456 -655 476 -654
rect 456 -658 476 -657
rect 456 -663 476 -662
rect 456 -666 476 -665
rect 14 -704 15 -684
rect 17 -704 18 -684
rect 22 -704 23 -684
rect 25 -704 26 -684
rect 44 -704 45 -684
rect 47 -704 48 -684
rect 52 -704 53 -684
rect 55 -704 56 -684
rect 84 -701 85 -681
rect 87 -701 88 -681
rect 107 -688 108 -668
rect 110 -688 111 -668
rect 147 -704 148 -684
rect 150 -704 151 -684
rect 248 -688 268 -687
rect 345 -687 346 -667
rect 348 -687 349 -667
rect 248 -691 268 -690
rect 248 -696 268 -695
rect 248 -699 268 -698
rect 457 -729 477 -728
rect 457 -732 477 -731
rect 457 -737 477 -736
rect 457 -740 477 -739
rect 457 -745 477 -744
rect 457 -748 477 -747
rect 457 -753 477 -752
rect 457 -756 477 -755
rect 464 -905 484 -904
rect 464 -908 484 -907
rect 464 -913 484 -912
rect 464 -916 484 -915
rect 458 -971 478 -970
rect 458 -974 478 -973
rect 458 -979 478 -978
rect 458 -982 478 -981
rect 458 -987 478 -986
rect 458 -990 478 -989
rect 14 -1052 15 -1032
rect 17 -1052 18 -1032
rect 22 -1052 23 -1032
rect 25 -1052 26 -1032
rect 44 -1052 45 -1032
rect 47 -1052 48 -1032
rect 52 -1052 53 -1032
rect 55 -1052 56 -1032
rect 84 -1049 85 -1029
rect 87 -1049 88 -1029
rect 107 -1036 108 -1016
rect 110 -1036 111 -1016
rect 147 -1052 148 -1032
rect 150 -1052 151 -1032
rect 262 -1038 263 -1018
rect 265 -1038 266 -1018
rect 285 -1038 286 -1018
rect 288 -1038 289 -1018
rect 238 -1075 239 -1055
rect 241 -1075 242 -1055
rect 458 -1053 478 -1052
rect 458 -1056 478 -1055
rect 458 -1061 478 -1060
rect 458 -1064 478 -1063
rect 458 -1069 478 -1068
rect 458 -1072 478 -1071
rect 458 -1077 478 -1076
rect 458 -1080 478 -1079
rect 465 -1140 479 -1139
rect 465 -1143 479 -1142
rect 465 -1148 479 -1147
rect 465 -1151 479 -1150
rect 12 -1193 13 -1173
rect 15 -1193 16 -1173
rect 20 -1193 21 -1173
rect 23 -1193 24 -1173
rect 42 -1193 43 -1173
rect 45 -1193 46 -1173
rect 50 -1193 51 -1173
rect 53 -1193 54 -1173
rect 82 -1190 83 -1170
rect 85 -1190 86 -1170
rect 105 -1177 106 -1157
rect 108 -1177 109 -1157
rect 344 -1172 345 -1152
rect 347 -1172 348 -1152
rect 465 -1156 479 -1155
rect 465 -1159 479 -1158
rect 465 -1164 479 -1163
rect 465 -1167 479 -1166
rect 145 -1193 146 -1173
rect 148 -1193 149 -1173
rect 246 -1177 266 -1176
rect 246 -1180 266 -1179
rect 246 -1185 266 -1184
rect 465 -1172 479 -1171
rect 465 -1175 479 -1174
rect 246 -1188 266 -1187
rect 464 -1224 478 -1223
rect 464 -1227 478 -1226
rect 464 -1232 478 -1231
rect 464 -1235 478 -1234
rect 464 -1240 478 -1239
rect 464 -1243 478 -1242
rect 464 -1248 478 -1247
rect 464 -1251 478 -1250
rect 464 -1256 478 -1255
rect 464 -1259 478 -1258
rect 463 -1400 483 -1399
rect 463 -1403 483 -1402
rect 463 -1408 483 -1407
rect 463 -1411 483 -1410
rect 457 -1466 477 -1465
rect 457 -1469 477 -1468
rect 457 -1474 477 -1473
rect 457 -1477 477 -1476
rect 457 -1482 477 -1481
rect 457 -1485 477 -1484
rect 12 -1542 13 -1522
rect 15 -1542 16 -1522
rect 20 -1542 21 -1522
rect 23 -1542 24 -1522
rect 42 -1542 43 -1522
rect 45 -1542 46 -1522
rect 50 -1542 51 -1522
rect 53 -1542 54 -1522
rect 82 -1539 83 -1519
rect 85 -1539 86 -1519
rect 105 -1526 106 -1506
rect 108 -1526 109 -1506
rect 145 -1542 146 -1522
rect 148 -1542 149 -1522
rect 261 -1528 262 -1508
rect 264 -1528 265 -1508
rect 284 -1528 285 -1508
rect 287 -1528 288 -1508
rect 237 -1565 238 -1545
rect 240 -1565 241 -1545
rect 457 -1548 477 -1547
rect 457 -1551 477 -1550
rect 457 -1556 477 -1555
rect 457 -1559 477 -1558
rect 457 -1564 477 -1563
rect 457 -1567 477 -1566
rect 457 -1572 477 -1571
rect 457 -1575 477 -1574
rect 464 -1635 478 -1634
rect 464 -1638 478 -1637
rect 12 -1683 13 -1663
rect 15 -1683 16 -1663
rect 20 -1683 21 -1663
rect 23 -1683 24 -1663
rect 42 -1683 43 -1663
rect 45 -1683 46 -1663
rect 50 -1683 51 -1663
rect 53 -1683 54 -1663
rect 82 -1680 83 -1660
rect 85 -1680 86 -1660
rect 105 -1667 106 -1647
rect 108 -1667 109 -1647
rect 344 -1658 345 -1638
rect 347 -1658 348 -1638
rect 464 -1643 478 -1642
rect 464 -1646 478 -1645
rect 464 -1651 478 -1650
rect 464 -1654 478 -1653
rect 145 -1683 146 -1663
rect 148 -1683 149 -1663
rect 245 -1667 265 -1666
rect 245 -1670 265 -1669
rect 245 -1675 265 -1674
rect 464 -1659 478 -1658
rect 464 -1662 478 -1661
rect 464 -1667 478 -1666
rect 464 -1670 478 -1669
rect 245 -1678 265 -1677
rect 454 -1739 474 -1738
rect 454 -1742 474 -1741
rect 454 -1747 474 -1746
rect 454 -1750 474 -1749
rect 454 -1755 474 -1754
rect 454 -1758 474 -1757
rect 454 -1763 474 -1762
rect 454 -1766 474 -1765
rect 454 -1771 474 -1770
rect 454 -1774 474 -1773
rect 454 -1779 474 -1778
rect 454 -1782 474 -1781
rect 451 -1832 471 -1831
rect 451 -1835 471 -1834
rect 451 -1840 471 -1839
rect 451 -1843 471 -1842
rect 451 -1848 471 -1847
rect 451 -1851 471 -1850
rect 451 -1856 471 -1855
rect 451 -1859 471 -1858
rect 451 -1864 471 -1863
rect 451 -1867 471 -1866
rect 451 -1872 471 -1871
rect 451 -1875 471 -1874
rect 12 -2012 13 -1992
rect 15 -2012 16 -1992
rect 20 -2012 21 -1992
rect 23 -2012 24 -1992
rect 42 -2012 43 -1992
rect 45 -2012 46 -1992
rect 50 -2012 51 -1992
rect 53 -2012 54 -1992
rect 82 -2009 83 -1989
rect 85 -2009 86 -1989
rect 105 -1996 106 -1976
rect 108 -1996 109 -1976
rect 145 -2012 146 -1992
rect 148 -2012 149 -1992
<< ndcontact >>
rect 12 23 16 33
rect 20 23 32 33
rect 42 23 46 33
rect 50 23 54 33
rect 58 23 62 33
rect 105 19 109 29
rect 113 19 117 29
rect 121 19 125 29
rect 145 22 149 32
rect 153 22 157 32
rect 260 40 264 50
rect 268 40 272 50
rect 283 34 287 44
rect 291 34 295 44
rect 490 45 510 49
rect 490 37 510 41
rect 490 29 510 33
rect 236 2 240 12
rect 244 2 248 12
rect 281 -75 301 -71
rect 490 -52 510 -48
rect 490 -60 510 -56
rect 490 -68 510 -64
rect 281 -83 301 -79
rect 281 -91 301 -87
rect 10 -115 14 -105
rect 18 -115 30 -105
rect 40 -115 44 -105
rect 48 -115 52 -105
rect 56 -115 60 -105
rect 338 -97 342 -87
rect 346 -97 350 -87
rect 103 -119 107 -109
rect 111 -119 115 -109
rect 119 -119 123 -109
rect 143 -116 147 -106
rect 151 -116 155 -106
rect 487 -216 507 -212
rect 487 -224 507 -220
rect 487 -232 507 -228
rect 10 -256 14 -246
rect 18 -256 30 -246
rect 40 -256 44 -246
rect 48 -256 52 -246
rect 56 -256 60 -246
rect 103 -260 107 -250
rect 111 -260 115 -250
rect 119 -260 123 -250
rect 143 -257 147 -247
rect 151 -257 155 -247
rect 260 -243 264 -233
rect 268 -243 272 -233
rect 283 -249 287 -239
rect 291 -249 295 -239
rect 236 -281 240 -271
rect 244 -281 248 -271
rect 481 -282 511 -278
rect 481 -290 511 -286
rect 481 -298 511 -294
rect 481 -306 511 -302
rect 281 -358 301 -354
rect 481 -357 511 -353
rect 281 -366 301 -362
rect 281 -374 301 -370
rect 481 -365 511 -361
rect 10 -398 14 -388
rect 18 -398 30 -388
rect 40 -398 44 -388
rect 48 -398 52 -388
rect 56 -398 60 -388
rect 341 -385 345 -375
rect 349 -385 353 -375
rect 481 -373 511 -369
rect 481 -381 511 -377
rect 103 -402 107 -392
rect 111 -402 115 -392
rect 119 -402 123 -392
rect 143 -399 147 -389
rect 151 -399 155 -389
rect 495 -490 515 -486
rect 495 -498 515 -494
rect 495 -506 515 -502
rect 489 -556 519 -552
rect 10 -585 14 -575
rect 18 -585 30 -575
rect 40 -585 44 -575
rect 48 -585 52 -575
rect 56 -585 60 -575
rect 103 -589 107 -579
rect 111 -589 115 -579
rect 119 -589 123 -579
rect 143 -586 147 -576
rect 151 -586 155 -576
rect 260 -572 264 -562
rect 268 -572 272 -562
rect 489 -564 519 -560
rect 283 -578 287 -568
rect 291 -578 295 -568
rect 489 -572 519 -568
rect 489 -580 519 -576
rect 236 -610 240 -600
rect 244 -610 248 -600
rect 489 -638 529 -634
rect 489 -646 529 -642
rect 489 -654 529 -650
rect 489 -662 529 -658
rect 281 -687 301 -683
rect 489 -670 529 -666
rect 281 -695 301 -691
rect 281 -703 301 -699
rect 10 -727 14 -717
rect 18 -727 30 -717
rect 40 -727 44 -717
rect 48 -727 52 -717
rect 56 -727 60 -717
rect 341 -711 345 -701
rect 349 -711 353 -701
rect 103 -731 107 -721
rect 111 -731 115 -721
rect 119 -731 123 -721
rect 143 -728 147 -718
rect 151 -728 155 -718
rect 490 -728 530 -724
rect 490 -736 530 -732
rect 490 -744 530 -740
rect 490 -752 530 -748
rect 490 -760 530 -756
rect 497 -904 517 -900
rect 497 -912 517 -908
rect 497 -920 517 -916
rect 491 -970 521 -966
rect 491 -978 521 -974
rect 491 -986 521 -982
rect 491 -994 521 -990
rect 10 -1075 14 -1065
rect 18 -1075 30 -1065
rect 40 -1075 44 -1065
rect 48 -1075 52 -1065
rect 56 -1075 60 -1065
rect 103 -1079 107 -1069
rect 111 -1079 115 -1069
rect 119 -1079 123 -1069
rect 143 -1076 147 -1066
rect 151 -1076 155 -1066
rect 258 -1061 262 -1051
rect 266 -1061 270 -1051
rect 491 -1052 531 -1048
rect 281 -1067 285 -1057
rect 289 -1067 293 -1057
rect 491 -1060 531 -1056
rect 491 -1068 531 -1064
rect 491 -1076 531 -1072
rect 491 -1084 531 -1080
rect 234 -1099 238 -1089
rect 242 -1099 246 -1089
rect 492 -1139 542 -1135
rect 492 -1147 542 -1143
rect 492 -1155 542 -1151
rect 492 -1163 542 -1159
rect 279 -1176 299 -1172
rect 279 -1184 299 -1180
rect 492 -1171 542 -1167
rect 492 -1179 542 -1175
rect 279 -1192 299 -1188
rect 8 -1216 12 -1206
rect 16 -1216 28 -1206
rect 38 -1216 42 -1206
rect 46 -1216 50 -1206
rect 54 -1216 58 -1206
rect 340 -1196 344 -1186
rect 348 -1196 352 -1186
rect 101 -1220 105 -1210
rect 109 -1220 113 -1210
rect 117 -1220 121 -1210
rect 141 -1217 145 -1207
rect 149 -1217 153 -1207
rect 491 -1223 541 -1219
rect 491 -1231 541 -1227
rect 491 -1239 541 -1235
rect 491 -1247 541 -1243
rect 491 -1255 541 -1251
rect 491 -1263 541 -1259
rect 496 -1399 516 -1395
rect 496 -1407 516 -1403
rect 496 -1415 516 -1411
rect 490 -1465 520 -1461
rect 490 -1473 520 -1469
rect 490 -1481 520 -1477
rect 490 -1489 520 -1485
rect 8 -1565 12 -1555
rect 16 -1565 28 -1555
rect 38 -1565 42 -1555
rect 46 -1565 50 -1555
rect 54 -1565 58 -1555
rect 101 -1569 105 -1559
rect 109 -1569 113 -1559
rect 117 -1569 121 -1559
rect 141 -1566 145 -1556
rect 149 -1566 153 -1556
rect 257 -1551 261 -1541
rect 265 -1551 269 -1541
rect 280 -1557 284 -1547
rect 288 -1557 292 -1547
rect 490 -1547 530 -1543
rect 490 -1555 530 -1551
rect 490 -1563 530 -1559
rect 490 -1571 530 -1567
rect 490 -1579 530 -1575
rect 233 -1589 237 -1579
rect 241 -1589 245 -1579
rect 491 -1634 541 -1630
rect 491 -1642 541 -1638
rect 491 -1650 541 -1646
rect 278 -1666 298 -1662
rect 278 -1674 298 -1670
rect 491 -1658 541 -1654
rect 491 -1666 541 -1662
rect 278 -1682 298 -1678
rect 340 -1682 344 -1672
rect 348 -1682 352 -1672
rect 491 -1674 541 -1670
rect 8 -1706 12 -1696
rect 16 -1706 28 -1696
rect 38 -1706 42 -1696
rect 46 -1706 50 -1696
rect 54 -1706 58 -1696
rect 101 -1710 105 -1700
rect 109 -1710 113 -1700
rect 117 -1710 121 -1700
rect 141 -1707 145 -1697
rect 149 -1707 153 -1697
rect 487 -1738 547 -1734
rect 487 -1746 547 -1742
rect 487 -1754 547 -1750
rect 487 -1762 547 -1758
rect 487 -1770 547 -1766
rect 487 -1778 547 -1774
rect 487 -1786 547 -1782
rect 484 -1831 544 -1827
rect 484 -1839 544 -1835
rect 484 -1847 544 -1843
rect 484 -1855 544 -1851
rect 484 -1863 544 -1859
rect 484 -1871 544 -1867
rect 484 -1879 544 -1875
rect 8 -2035 12 -2025
rect 16 -2035 28 -2025
rect 38 -2035 42 -2025
rect 46 -2035 50 -2025
rect 54 -2035 58 -2025
rect 101 -2039 105 -2029
rect 109 -2039 113 -2029
rect 117 -2039 121 -2029
rect 141 -2036 145 -2026
rect 149 -2036 153 -2026
<< pdcontact >>
rect 12 46 16 66
rect 20 46 24 66
rect 28 46 32 66
rect 42 46 46 66
rect 50 46 54 66
rect 58 46 62 66
rect 82 49 86 69
rect 90 49 94 69
rect 105 62 109 82
rect 113 62 125 82
rect 145 46 149 66
rect 153 46 157 66
rect 260 63 264 83
rect 268 63 272 83
rect 283 63 287 83
rect 291 63 295 83
rect 236 26 240 46
rect 244 26 248 46
rect 457 45 477 49
rect 457 37 477 41
rect 457 29 477 33
rect 10 -92 14 -72
rect 18 -92 22 -72
rect 26 -92 30 -72
rect 40 -92 44 -72
rect 48 -92 52 -72
rect 56 -92 60 -72
rect 80 -89 84 -69
rect 88 -89 92 -69
rect 103 -76 107 -56
rect 111 -76 123 -56
rect 143 -92 147 -72
rect 151 -92 155 -72
rect 248 -75 268 -71
rect 338 -73 342 -53
rect 346 -73 350 -53
rect 457 -52 477 -48
rect 457 -60 477 -56
rect 457 -68 477 -64
rect 248 -83 268 -79
rect 248 -91 268 -87
rect 10 -233 14 -213
rect 18 -233 22 -213
rect 26 -233 30 -213
rect 40 -233 44 -213
rect 48 -233 52 -213
rect 56 -233 60 -213
rect 80 -230 84 -210
rect 88 -230 92 -210
rect 103 -217 107 -197
rect 111 -217 123 -197
rect 143 -233 147 -213
rect 151 -233 155 -213
rect 260 -220 264 -200
rect 268 -220 272 -200
rect 283 -220 287 -200
rect 291 -220 295 -200
rect 454 -216 474 -212
rect 454 -224 474 -220
rect 454 -232 474 -228
rect 236 -257 240 -237
rect 244 -257 248 -237
rect 448 -282 468 -278
rect 448 -290 468 -286
rect 448 -298 468 -294
rect 448 -306 468 -302
rect 10 -375 14 -355
rect 18 -375 22 -355
rect 26 -375 30 -355
rect 40 -375 44 -355
rect 48 -375 52 -355
rect 56 -375 60 -355
rect 80 -372 84 -352
rect 88 -372 92 -352
rect 103 -359 107 -339
rect 111 -359 123 -339
rect 143 -375 147 -355
rect 151 -375 155 -355
rect 248 -358 268 -354
rect 341 -361 345 -341
rect 349 -361 353 -341
rect 448 -357 468 -353
rect 248 -366 268 -362
rect 248 -374 268 -370
rect 448 -365 468 -361
rect 448 -373 468 -369
rect 448 -381 468 -377
rect 462 -490 482 -486
rect 462 -498 482 -494
rect 462 -506 482 -502
rect 10 -562 14 -542
rect 18 -562 22 -542
rect 26 -562 30 -542
rect 40 -562 44 -542
rect 48 -562 52 -542
rect 56 -562 60 -542
rect 80 -559 84 -539
rect 88 -559 92 -539
rect 103 -546 107 -526
rect 111 -546 123 -526
rect 143 -562 147 -542
rect 151 -562 155 -542
rect 260 -549 264 -529
rect 268 -549 272 -529
rect 283 -549 287 -529
rect 291 -549 295 -529
rect 456 -556 476 -552
rect 236 -586 240 -566
rect 244 -586 248 -566
rect 456 -564 476 -560
rect 456 -572 476 -568
rect 456 -580 476 -576
rect 456 -638 476 -634
rect 456 -646 476 -642
rect 456 -654 476 -650
rect 456 -662 476 -658
rect 10 -704 14 -684
rect 18 -704 22 -684
rect 26 -704 30 -684
rect 40 -704 44 -684
rect 48 -704 52 -684
rect 56 -704 60 -684
rect 80 -701 84 -681
rect 88 -701 92 -681
rect 103 -688 107 -668
rect 111 -688 123 -668
rect 143 -704 147 -684
rect 151 -704 155 -684
rect 248 -687 268 -683
rect 341 -687 345 -667
rect 349 -687 353 -667
rect 456 -670 476 -666
rect 248 -695 268 -691
rect 248 -703 268 -699
rect 457 -728 477 -724
rect 457 -736 477 -732
rect 457 -744 477 -740
rect 457 -752 477 -748
rect 457 -760 477 -756
rect 464 -904 484 -900
rect 464 -912 484 -908
rect 464 -920 484 -916
rect 458 -970 478 -966
rect 458 -978 478 -974
rect 458 -986 478 -982
rect 458 -994 478 -990
rect 10 -1052 14 -1032
rect 18 -1052 22 -1032
rect 26 -1052 30 -1032
rect 40 -1052 44 -1032
rect 48 -1052 52 -1032
rect 56 -1052 60 -1032
rect 80 -1049 84 -1029
rect 88 -1049 92 -1029
rect 103 -1036 107 -1016
rect 111 -1036 123 -1016
rect 143 -1052 147 -1032
rect 151 -1052 155 -1032
rect 258 -1038 262 -1018
rect 266 -1038 270 -1018
rect 281 -1038 285 -1018
rect 289 -1038 293 -1018
rect 234 -1075 238 -1055
rect 242 -1075 246 -1055
rect 458 -1052 478 -1048
rect 458 -1060 478 -1056
rect 458 -1068 478 -1064
rect 458 -1076 478 -1072
rect 458 -1084 478 -1080
rect 465 -1139 479 -1135
rect 465 -1147 479 -1143
rect 8 -1193 12 -1173
rect 16 -1193 20 -1173
rect 24 -1193 28 -1173
rect 38 -1193 42 -1173
rect 46 -1193 50 -1173
rect 54 -1193 58 -1173
rect 78 -1190 82 -1170
rect 86 -1190 90 -1170
rect 101 -1177 105 -1157
rect 109 -1177 121 -1157
rect 340 -1172 344 -1152
rect 348 -1172 352 -1152
rect 465 -1155 479 -1151
rect 465 -1163 479 -1159
rect 465 -1171 479 -1167
rect 141 -1193 145 -1173
rect 149 -1193 153 -1173
rect 246 -1176 266 -1172
rect 246 -1184 266 -1180
rect 465 -1179 479 -1175
rect 246 -1192 266 -1188
rect 464 -1223 478 -1219
rect 464 -1231 478 -1227
rect 464 -1239 478 -1235
rect 464 -1247 478 -1243
rect 464 -1255 478 -1251
rect 464 -1263 478 -1259
rect 463 -1399 483 -1395
rect 463 -1407 483 -1403
rect 463 -1415 483 -1411
rect 457 -1465 477 -1461
rect 457 -1473 477 -1469
rect 457 -1481 477 -1477
rect 457 -1489 477 -1485
rect 8 -1542 12 -1522
rect 16 -1542 20 -1522
rect 24 -1542 28 -1522
rect 38 -1542 42 -1522
rect 46 -1542 50 -1522
rect 54 -1542 58 -1522
rect 78 -1539 82 -1519
rect 86 -1539 90 -1519
rect 101 -1526 105 -1506
rect 109 -1526 121 -1506
rect 141 -1542 145 -1522
rect 149 -1542 153 -1522
rect 257 -1528 261 -1508
rect 265 -1528 269 -1508
rect 280 -1528 284 -1508
rect 288 -1528 292 -1508
rect 233 -1565 237 -1545
rect 241 -1565 245 -1545
rect 457 -1547 477 -1543
rect 457 -1555 477 -1551
rect 457 -1563 477 -1559
rect 457 -1571 477 -1567
rect 457 -1579 477 -1575
rect 464 -1634 478 -1630
rect 8 -1683 12 -1663
rect 16 -1683 20 -1663
rect 24 -1683 28 -1663
rect 38 -1683 42 -1663
rect 46 -1683 50 -1663
rect 54 -1683 58 -1663
rect 78 -1680 82 -1660
rect 86 -1680 90 -1660
rect 101 -1667 105 -1647
rect 109 -1667 121 -1647
rect 340 -1658 344 -1638
rect 348 -1658 352 -1638
rect 464 -1642 478 -1638
rect 464 -1650 478 -1646
rect 464 -1658 478 -1654
rect 141 -1683 145 -1663
rect 149 -1683 153 -1663
rect 245 -1666 265 -1662
rect 245 -1674 265 -1670
rect 464 -1666 478 -1662
rect 245 -1682 265 -1678
rect 464 -1674 478 -1670
rect 454 -1738 474 -1734
rect 454 -1746 474 -1742
rect 454 -1754 474 -1750
rect 454 -1762 474 -1758
rect 454 -1770 474 -1766
rect 454 -1778 474 -1774
rect 454 -1786 474 -1782
rect 451 -1831 471 -1827
rect 451 -1839 471 -1835
rect 451 -1847 471 -1843
rect 451 -1855 471 -1851
rect 451 -1863 471 -1859
rect 451 -1871 471 -1867
rect 451 -1879 471 -1875
rect 8 -2012 12 -1992
rect 16 -2012 20 -1992
rect 24 -2012 28 -1992
rect 38 -2012 42 -1992
rect 46 -2012 50 -1992
rect 54 -2012 58 -1992
rect 78 -2009 82 -1989
rect 86 -2009 90 -1989
rect 101 -1996 105 -1976
rect 109 -1996 121 -1976
rect 141 -2012 145 -1992
rect 149 -2012 153 -1992
<< psubstratepcontact >>
rect 514 29 518 33
rect 0 0 4 5
rect 236 -6 240 -2
rect 514 -68 518 -64
rect 305 -91 309 -87
rect 338 -105 342 -101
rect -2 -138 2 -133
rect 511 -232 515 -228
rect -2 -279 2 -274
rect 236 -289 240 -285
rect 516 -306 520 -302
rect 305 -374 309 -370
rect 516 -381 520 -377
rect 341 -393 345 -389
rect -2 -421 2 -416
rect 519 -506 523 -502
rect 524 -580 528 -576
rect -2 -608 2 -603
rect 236 -618 240 -614
rect 534 -670 538 -666
rect 305 -703 309 -699
rect 341 -719 345 -715
rect -2 -750 2 -745
rect 535 -760 539 -756
rect 521 -920 525 -916
rect 526 -994 530 -990
rect 536 -1084 540 -1080
rect -2 -1098 2 -1093
rect 234 -1107 238 -1103
rect 549 -1179 553 -1175
rect 303 -1192 307 -1188
rect 340 -1204 344 -1200
rect -4 -1239 0 -1234
rect 548 -1263 552 -1259
rect 520 -1415 524 -1411
rect 525 -1489 529 -1485
rect 535 -1579 539 -1575
rect -4 -1588 0 -1583
rect 233 -1597 237 -1593
rect 302 -1682 306 -1678
rect 548 -1674 552 -1670
rect 340 -1690 344 -1686
rect -4 -1729 0 -1724
rect 552 -1786 556 -1782
rect 549 -1879 553 -1875
rect -4 -2058 0 -2053
<< nsubstratencontact >>
rect 155 90 159 94
rect 236 50 240 54
rect 448 29 452 33
rect 153 -48 157 -44
rect 338 -49 342 -45
rect 448 -68 452 -64
rect 239 -91 243 -87
rect 153 -189 157 -185
rect 236 -233 240 -229
rect 445 -232 449 -228
rect 439 -306 443 -302
rect 153 -331 157 -327
rect 341 -337 345 -333
rect 239 -374 243 -370
rect 439 -381 443 -377
rect 453 -506 457 -502
rect 153 -518 157 -514
rect 236 -562 240 -558
rect 447 -580 451 -576
rect 153 -660 157 -656
rect 341 -663 345 -659
rect 447 -670 451 -666
rect 239 -703 243 -699
rect 448 -760 452 -756
rect 455 -920 459 -916
rect 449 -994 453 -990
rect 153 -1008 157 -1004
rect 234 -1051 238 -1047
rect 449 -1084 453 -1080
rect 151 -1149 155 -1145
rect 340 -1148 344 -1144
rect 452 -1179 456 -1175
rect 237 -1192 241 -1188
rect 451 -1263 455 -1259
rect 454 -1415 458 -1411
rect 448 -1489 452 -1485
rect 151 -1498 155 -1494
rect 233 -1541 237 -1537
rect 448 -1579 452 -1575
rect 340 -1634 344 -1630
rect 151 -1639 155 -1635
rect 236 -1682 240 -1678
rect 451 -1674 455 -1670
rect 445 -1786 449 -1782
rect 442 -1879 446 -1875
rect 151 -1968 155 -1964
<< polysilicon >>
rect 110 82 112 86
rect 265 83 267 96
rect 288 83 290 87
rect 17 66 19 70
rect 25 66 27 70
rect 47 66 49 70
rect 55 66 57 70
rect 87 69 89 73
rect 150 66 152 70
rect 17 33 19 46
rect 25 42 27 46
rect 47 33 49 46
rect 55 33 57 46
rect 87 45 89 49
rect 110 43 112 62
rect 265 50 267 63
rect 288 59 290 63
rect 241 46 243 49
rect 110 29 112 34
rect 118 29 120 33
rect 150 32 152 46
rect 17 19 19 23
rect 47 19 49 23
rect 55 19 57 23
rect 288 44 290 51
rect 265 37 267 40
rect 440 42 457 44
rect 477 42 490 44
rect 510 42 513 44
rect 440 34 457 36
rect 477 34 490 36
rect 510 34 513 36
rect 288 31 290 34
rect 150 19 152 22
rect 110 15 112 19
rect 118 15 120 19
rect 241 12 243 26
rect 241 -1 243 2
rect 108 -56 110 -52
rect 343 -53 345 -50
rect 15 -72 17 -68
rect 23 -72 25 -68
rect 45 -72 47 -68
rect 53 -72 55 -68
rect 85 -69 87 -65
rect 148 -72 150 -68
rect 15 -105 17 -92
rect 23 -96 25 -92
rect 45 -105 47 -92
rect 53 -105 55 -92
rect 85 -93 87 -89
rect 108 -95 110 -76
rect 440 -55 457 -53
rect 477 -55 490 -53
rect 510 -55 513 -53
rect 440 -63 457 -61
rect 477 -63 490 -61
rect 510 -63 513 -61
rect 231 -78 248 -76
rect 268 -78 281 -76
rect 301 -78 304 -76
rect 231 -86 248 -84
rect 268 -86 281 -84
rect 301 -86 304 -84
rect 343 -87 345 -73
rect 108 -109 110 -104
rect 116 -109 118 -105
rect 148 -106 150 -92
rect 343 -100 345 -97
rect 15 -119 17 -115
rect 45 -119 47 -115
rect 53 -119 55 -115
rect 148 -119 150 -116
rect 108 -123 110 -119
rect 116 -123 118 -119
rect 108 -197 110 -193
rect 15 -213 17 -209
rect 23 -213 25 -209
rect 45 -213 47 -209
rect 53 -213 55 -209
rect 85 -210 87 -206
rect 265 -200 267 -187
rect 288 -200 290 -196
rect 148 -213 150 -209
rect 15 -246 17 -233
rect 23 -237 25 -233
rect 45 -246 47 -233
rect 53 -246 55 -233
rect 85 -234 87 -230
rect 108 -236 110 -217
rect 437 -219 454 -217
rect 474 -219 487 -217
rect 507 -219 510 -217
rect 265 -233 267 -220
rect 288 -224 290 -220
rect 437 -227 454 -225
rect 474 -227 487 -225
rect 507 -227 510 -225
rect 108 -250 110 -245
rect 116 -250 118 -246
rect 148 -247 150 -233
rect 241 -237 243 -234
rect 15 -260 17 -256
rect 45 -260 47 -256
rect 53 -260 55 -256
rect 288 -239 290 -232
rect 265 -246 267 -243
rect 288 -252 290 -249
rect 148 -260 150 -257
rect 108 -264 110 -260
rect 116 -264 118 -260
rect 241 -271 243 -257
rect 241 -284 243 -281
rect 431 -285 448 -283
rect 468 -285 481 -283
rect 511 -285 514 -283
rect 431 -293 448 -291
rect 468 -293 481 -291
rect 511 -293 514 -291
rect 431 -301 448 -299
rect 468 -301 481 -299
rect 511 -301 514 -299
rect 108 -339 110 -335
rect 15 -355 17 -351
rect 23 -355 25 -351
rect 45 -355 47 -351
rect 53 -355 55 -351
rect 85 -352 87 -348
rect 346 -341 348 -338
rect 148 -355 150 -351
rect 15 -388 17 -375
rect 23 -379 25 -375
rect 45 -388 47 -375
rect 53 -388 55 -375
rect 85 -376 87 -372
rect 108 -378 110 -359
rect 231 -361 248 -359
rect 268 -361 281 -359
rect 301 -361 304 -359
rect 431 -360 448 -358
rect 468 -360 481 -358
rect 511 -360 514 -358
rect 231 -369 248 -367
rect 268 -369 281 -367
rect 301 -369 304 -367
rect 346 -375 348 -361
rect 431 -368 448 -366
rect 468 -368 481 -366
rect 511 -368 514 -366
rect 108 -392 110 -387
rect 116 -392 118 -388
rect 148 -389 150 -375
rect 431 -376 448 -374
rect 468 -376 481 -374
rect 511 -376 514 -374
rect 346 -388 348 -385
rect 15 -402 17 -398
rect 45 -402 47 -398
rect 53 -402 55 -398
rect 148 -402 150 -399
rect 108 -406 110 -402
rect 116 -406 118 -402
rect 445 -493 462 -491
rect 482 -493 495 -491
rect 515 -493 518 -491
rect 445 -501 462 -499
rect 482 -501 495 -499
rect 515 -501 518 -499
rect 108 -526 110 -522
rect 15 -542 17 -538
rect 23 -542 25 -538
rect 45 -542 47 -538
rect 53 -542 55 -538
rect 85 -539 87 -535
rect 265 -529 267 -516
rect 288 -529 290 -525
rect 148 -542 150 -538
rect 15 -575 17 -562
rect 23 -566 25 -562
rect 45 -575 47 -562
rect 53 -575 55 -562
rect 85 -563 87 -559
rect 108 -565 110 -546
rect 265 -562 267 -549
rect 288 -553 290 -549
rect 439 -559 456 -557
rect 476 -559 489 -557
rect 519 -559 522 -557
rect 108 -579 110 -574
rect 116 -579 118 -575
rect 148 -576 150 -562
rect 241 -566 243 -563
rect 15 -589 17 -585
rect 45 -589 47 -585
rect 53 -589 55 -585
rect 288 -568 290 -561
rect 439 -567 456 -565
rect 476 -567 489 -565
rect 519 -567 522 -565
rect 265 -575 267 -572
rect 439 -575 456 -573
rect 476 -575 489 -573
rect 519 -575 522 -573
rect 288 -581 290 -578
rect 148 -589 150 -586
rect 108 -593 110 -589
rect 116 -593 118 -589
rect 241 -600 243 -586
rect 241 -613 243 -610
rect 439 -641 456 -639
rect 476 -641 489 -639
rect 529 -641 532 -639
rect 439 -649 456 -647
rect 476 -649 489 -647
rect 529 -649 532 -647
rect 439 -657 456 -655
rect 476 -657 489 -655
rect 529 -657 532 -655
rect 108 -668 110 -664
rect 346 -667 348 -664
rect 439 -665 456 -663
rect 476 -665 489 -663
rect 529 -665 532 -663
rect 15 -684 17 -680
rect 23 -684 25 -680
rect 45 -684 47 -680
rect 53 -684 55 -680
rect 85 -681 87 -677
rect 148 -684 150 -680
rect 15 -717 17 -704
rect 23 -708 25 -704
rect 45 -717 47 -704
rect 53 -717 55 -704
rect 85 -705 87 -701
rect 108 -707 110 -688
rect 231 -690 248 -688
rect 268 -690 281 -688
rect 301 -690 304 -688
rect 231 -698 248 -696
rect 268 -698 281 -696
rect 301 -698 304 -696
rect 346 -701 348 -687
rect 108 -721 110 -716
rect 116 -721 118 -717
rect 148 -718 150 -704
rect 346 -714 348 -711
rect 15 -731 17 -727
rect 45 -731 47 -727
rect 53 -731 55 -727
rect 148 -731 150 -728
rect 440 -731 457 -729
rect 477 -731 490 -729
rect 530 -731 533 -729
rect 108 -735 110 -731
rect 116 -735 118 -731
rect 440 -739 457 -737
rect 477 -739 490 -737
rect 530 -739 533 -737
rect 440 -747 457 -745
rect 477 -747 490 -745
rect 530 -747 533 -745
rect 440 -755 457 -753
rect 477 -755 490 -753
rect 530 -755 533 -753
rect 447 -907 464 -905
rect 484 -907 497 -905
rect 517 -907 520 -905
rect 447 -915 464 -913
rect 484 -915 497 -913
rect 517 -915 520 -913
rect 441 -973 458 -971
rect 478 -973 491 -971
rect 521 -973 524 -971
rect 441 -981 458 -979
rect 478 -981 491 -979
rect 521 -981 524 -979
rect 441 -989 458 -987
rect 478 -989 491 -987
rect 521 -989 524 -987
rect 108 -1016 110 -1012
rect 15 -1032 17 -1028
rect 23 -1032 25 -1028
rect 45 -1032 47 -1028
rect 53 -1032 55 -1028
rect 85 -1029 87 -1025
rect 263 -1018 265 -1005
rect 286 -1018 288 -1014
rect 148 -1032 150 -1028
rect 15 -1065 17 -1052
rect 23 -1056 25 -1052
rect 45 -1065 47 -1052
rect 53 -1065 55 -1052
rect 85 -1053 87 -1049
rect 108 -1055 110 -1036
rect 263 -1051 265 -1038
rect 286 -1042 288 -1038
rect 108 -1069 110 -1064
rect 116 -1069 118 -1065
rect 148 -1066 150 -1052
rect 239 -1055 241 -1052
rect 15 -1079 17 -1075
rect 45 -1079 47 -1075
rect 53 -1079 55 -1075
rect 286 -1057 288 -1050
rect 441 -1055 458 -1053
rect 478 -1055 491 -1053
rect 531 -1055 534 -1053
rect 263 -1064 265 -1061
rect 441 -1063 458 -1061
rect 478 -1063 491 -1061
rect 531 -1063 534 -1061
rect 286 -1070 288 -1067
rect 441 -1071 458 -1069
rect 478 -1071 491 -1069
rect 531 -1071 534 -1069
rect 148 -1079 150 -1076
rect 108 -1083 110 -1079
rect 116 -1083 118 -1079
rect 239 -1089 241 -1075
rect 441 -1079 458 -1077
rect 478 -1079 491 -1077
rect 531 -1079 534 -1077
rect 239 -1102 241 -1099
rect 442 -1142 465 -1140
rect 479 -1142 492 -1140
rect 542 -1142 545 -1140
rect 345 -1152 347 -1149
rect 442 -1150 465 -1148
rect 479 -1150 492 -1148
rect 542 -1150 545 -1148
rect 106 -1157 108 -1153
rect 13 -1173 15 -1169
rect 21 -1173 23 -1169
rect 43 -1173 45 -1169
rect 51 -1173 53 -1169
rect 83 -1170 85 -1166
rect 146 -1173 148 -1169
rect 442 -1158 465 -1156
rect 479 -1158 492 -1156
rect 542 -1158 545 -1156
rect 442 -1166 465 -1164
rect 479 -1166 492 -1164
rect 542 -1166 545 -1164
rect 13 -1206 15 -1193
rect 21 -1197 23 -1193
rect 43 -1206 45 -1193
rect 51 -1206 53 -1193
rect 83 -1194 85 -1190
rect 106 -1196 108 -1177
rect 229 -1179 246 -1177
rect 266 -1179 279 -1177
rect 299 -1179 302 -1177
rect 229 -1187 246 -1185
rect 266 -1187 279 -1185
rect 299 -1187 302 -1185
rect 345 -1186 347 -1172
rect 442 -1174 465 -1172
rect 479 -1174 492 -1172
rect 542 -1174 545 -1172
rect 106 -1210 108 -1205
rect 114 -1210 116 -1206
rect 146 -1207 148 -1193
rect 345 -1199 347 -1196
rect 13 -1220 15 -1216
rect 43 -1220 45 -1216
rect 51 -1220 53 -1216
rect 146 -1220 148 -1217
rect 106 -1224 108 -1220
rect 114 -1224 116 -1220
rect 441 -1226 464 -1224
rect 478 -1226 491 -1224
rect 541 -1226 544 -1224
rect 441 -1234 464 -1232
rect 478 -1234 491 -1232
rect 541 -1234 544 -1232
rect 441 -1242 464 -1240
rect 478 -1242 491 -1240
rect 541 -1242 544 -1240
rect 441 -1250 464 -1248
rect 478 -1250 491 -1248
rect 541 -1250 544 -1248
rect 441 -1258 464 -1256
rect 478 -1258 491 -1256
rect 541 -1258 544 -1256
rect 446 -1402 463 -1400
rect 483 -1402 496 -1400
rect 516 -1402 519 -1400
rect 446 -1410 463 -1408
rect 483 -1410 496 -1408
rect 516 -1410 519 -1408
rect 440 -1468 457 -1466
rect 477 -1468 490 -1466
rect 520 -1468 523 -1466
rect 440 -1476 457 -1474
rect 477 -1476 490 -1474
rect 520 -1476 523 -1474
rect 440 -1484 457 -1482
rect 477 -1484 490 -1482
rect 520 -1484 523 -1482
rect 106 -1506 108 -1502
rect 13 -1522 15 -1518
rect 21 -1522 23 -1518
rect 43 -1522 45 -1518
rect 51 -1522 53 -1518
rect 83 -1519 85 -1515
rect 262 -1508 264 -1495
rect 285 -1508 287 -1504
rect 146 -1522 148 -1518
rect 13 -1555 15 -1542
rect 21 -1546 23 -1542
rect 43 -1555 45 -1542
rect 51 -1555 53 -1542
rect 83 -1543 85 -1539
rect 106 -1545 108 -1526
rect 262 -1541 264 -1528
rect 285 -1532 287 -1528
rect 106 -1559 108 -1554
rect 114 -1559 116 -1555
rect 146 -1556 148 -1542
rect 238 -1545 240 -1542
rect 13 -1569 15 -1565
rect 43 -1569 45 -1565
rect 51 -1569 53 -1565
rect 285 -1547 287 -1540
rect 262 -1554 264 -1551
rect 440 -1550 457 -1548
rect 477 -1550 490 -1548
rect 530 -1550 533 -1548
rect 285 -1560 287 -1557
rect 440 -1558 457 -1556
rect 477 -1558 490 -1556
rect 530 -1558 533 -1556
rect 146 -1569 148 -1566
rect 106 -1573 108 -1569
rect 114 -1573 116 -1569
rect 238 -1579 240 -1565
rect 440 -1566 457 -1564
rect 477 -1566 490 -1564
rect 530 -1566 533 -1564
rect 440 -1574 457 -1572
rect 477 -1574 490 -1572
rect 530 -1574 533 -1572
rect 238 -1592 240 -1589
rect 345 -1638 347 -1635
rect 441 -1637 464 -1635
rect 478 -1637 491 -1635
rect 541 -1637 544 -1635
rect 106 -1647 108 -1643
rect 13 -1663 15 -1659
rect 21 -1663 23 -1659
rect 43 -1663 45 -1659
rect 51 -1663 53 -1659
rect 83 -1660 85 -1656
rect 441 -1645 464 -1643
rect 478 -1645 491 -1643
rect 541 -1645 544 -1643
rect 441 -1653 464 -1651
rect 478 -1653 491 -1651
rect 541 -1653 544 -1651
rect 146 -1663 148 -1659
rect 13 -1696 15 -1683
rect 21 -1687 23 -1683
rect 43 -1696 45 -1683
rect 51 -1696 53 -1683
rect 83 -1684 85 -1680
rect 106 -1686 108 -1667
rect 228 -1669 245 -1667
rect 265 -1669 278 -1667
rect 298 -1669 301 -1667
rect 345 -1672 347 -1658
rect 441 -1661 464 -1659
rect 478 -1661 491 -1659
rect 541 -1661 544 -1659
rect 441 -1669 464 -1667
rect 478 -1669 491 -1667
rect 541 -1669 544 -1667
rect 228 -1677 245 -1675
rect 265 -1677 278 -1675
rect 298 -1677 301 -1675
rect 106 -1700 108 -1695
rect 114 -1700 116 -1696
rect 146 -1697 148 -1683
rect 345 -1685 347 -1682
rect 13 -1710 15 -1706
rect 43 -1710 45 -1706
rect 51 -1710 53 -1706
rect 146 -1710 148 -1707
rect 106 -1714 108 -1710
rect 114 -1714 116 -1710
rect 437 -1741 454 -1739
rect 474 -1741 487 -1739
rect 547 -1741 550 -1739
rect 437 -1749 454 -1747
rect 474 -1749 487 -1747
rect 547 -1749 550 -1747
rect 437 -1757 454 -1755
rect 474 -1757 487 -1755
rect 547 -1757 550 -1755
rect 437 -1765 454 -1763
rect 474 -1765 487 -1763
rect 547 -1765 550 -1763
rect 437 -1773 454 -1771
rect 474 -1773 487 -1771
rect 547 -1773 550 -1771
rect 437 -1781 454 -1779
rect 474 -1781 487 -1779
rect 547 -1781 550 -1779
rect 434 -1834 451 -1832
rect 471 -1834 484 -1832
rect 544 -1834 547 -1832
rect 434 -1842 451 -1840
rect 471 -1842 484 -1840
rect 544 -1842 547 -1840
rect 434 -1850 451 -1848
rect 471 -1850 484 -1848
rect 544 -1850 547 -1848
rect 434 -1858 451 -1856
rect 471 -1858 484 -1856
rect 544 -1858 547 -1856
rect 434 -1866 451 -1864
rect 471 -1866 484 -1864
rect 544 -1866 547 -1864
rect 434 -1874 451 -1872
rect 471 -1874 484 -1872
rect 544 -1874 547 -1872
rect 106 -1976 108 -1972
rect 13 -1992 15 -1988
rect 21 -1992 23 -1988
rect 43 -1992 45 -1988
rect 51 -1992 53 -1988
rect 83 -1989 85 -1985
rect 146 -1992 148 -1988
rect 13 -2025 15 -2012
rect 21 -2016 23 -2012
rect 43 -2025 45 -2012
rect 51 -2025 53 -2012
rect 83 -2013 85 -2009
rect 106 -2015 108 -1996
rect 106 -2029 108 -2024
rect 114 -2029 116 -2025
rect 146 -2026 148 -2012
rect 13 -2039 15 -2035
rect 43 -2039 45 -2035
rect 51 -2039 53 -2035
rect 146 -2039 148 -2036
rect 106 -2043 108 -2039
rect 114 -2043 116 -2039
<< polycontact >>
rect 265 96 269 100
rect 285 87 290 92
rect 17 70 21 74
rect 54 70 58 74
rect 87 73 91 77
rect 106 55 110 59
rect 106 43 110 47
rect 106 32 110 36
rect 146 35 150 39
rect 436 42 440 46
rect 436 34 440 38
rect 288 27 292 31
rect 237 15 241 19
rect 15 -68 19 -64
rect 52 -68 56 -64
rect 85 -65 89 -61
rect 104 -83 108 -79
rect 104 -95 108 -91
rect 227 -78 231 -74
rect 436 -55 440 -51
rect 436 -63 440 -59
rect 227 -86 231 -82
rect 339 -84 343 -80
rect 104 -106 108 -102
rect 144 -103 148 -99
rect 265 -187 269 -183
rect 15 -209 19 -205
rect 52 -209 56 -205
rect 85 -206 89 -202
rect 285 -196 290 -191
rect 104 -224 108 -220
rect 104 -236 108 -232
rect 433 -219 437 -215
rect 433 -227 437 -223
rect 104 -247 108 -243
rect 144 -244 148 -240
rect 288 -256 292 -252
rect 237 -268 241 -264
rect 427 -285 431 -281
rect 427 -293 431 -289
rect 427 -301 431 -297
rect 15 -351 19 -347
rect 52 -351 56 -347
rect 85 -348 89 -344
rect 104 -366 108 -362
rect 104 -378 108 -374
rect 227 -361 231 -357
rect 427 -360 431 -356
rect 227 -369 231 -365
rect 342 -372 346 -368
rect 427 -368 431 -364
rect 104 -389 108 -385
rect 144 -386 148 -382
rect 427 -376 431 -372
rect 441 -493 445 -489
rect 441 -501 445 -497
rect 265 -516 269 -512
rect 15 -538 19 -534
rect 52 -538 56 -534
rect 85 -535 89 -531
rect 285 -525 290 -520
rect 104 -553 108 -549
rect 104 -565 108 -561
rect 435 -559 439 -555
rect 104 -576 108 -572
rect 144 -573 148 -569
rect 435 -567 439 -563
rect 435 -575 439 -571
rect 288 -585 292 -581
rect 237 -597 241 -593
rect 435 -641 439 -637
rect 435 -649 439 -645
rect 435 -657 439 -653
rect 435 -665 439 -661
rect 15 -680 19 -676
rect 52 -680 56 -676
rect 85 -677 89 -673
rect 104 -695 108 -691
rect 104 -707 108 -703
rect 227 -690 231 -686
rect 227 -698 231 -694
rect 342 -698 346 -694
rect 104 -718 108 -714
rect 144 -715 148 -711
rect 436 -731 440 -727
rect 436 -739 440 -735
rect 436 -747 440 -743
rect 436 -755 440 -751
rect 443 -907 447 -903
rect 443 -915 447 -911
rect 437 -973 441 -969
rect 437 -981 441 -977
rect 437 -989 441 -985
rect 263 -1005 267 -1001
rect 15 -1028 19 -1024
rect 52 -1028 56 -1024
rect 85 -1025 89 -1021
rect 283 -1014 288 -1009
rect 104 -1043 108 -1039
rect 104 -1055 108 -1051
rect 104 -1066 108 -1062
rect 144 -1063 148 -1059
rect 437 -1055 441 -1051
rect 437 -1063 441 -1059
rect 286 -1074 290 -1070
rect 437 -1071 441 -1067
rect 235 -1086 239 -1082
rect 437 -1079 441 -1075
rect 438 -1143 442 -1139
rect 438 -1151 442 -1147
rect 13 -1169 17 -1165
rect 50 -1169 54 -1165
rect 83 -1166 87 -1162
rect 438 -1159 442 -1155
rect 438 -1167 442 -1163
rect 102 -1184 106 -1180
rect 102 -1196 106 -1192
rect 225 -1179 229 -1175
rect 225 -1187 229 -1183
rect 341 -1183 345 -1179
rect 438 -1175 442 -1171
rect 102 -1207 106 -1203
rect 142 -1204 146 -1200
rect 437 -1227 441 -1223
rect 437 -1235 441 -1231
rect 437 -1243 441 -1239
rect 437 -1251 441 -1247
rect 437 -1259 441 -1255
rect 442 -1402 446 -1398
rect 442 -1410 446 -1406
rect 436 -1468 440 -1464
rect 436 -1476 440 -1472
rect 436 -1484 440 -1480
rect 262 -1495 266 -1491
rect 13 -1518 17 -1514
rect 50 -1518 54 -1514
rect 83 -1515 87 -1511
rect 282 -1504 287 -1499
rect 102 -1533 106 -1529
rect 102 -1545 106 -1541
rect 102 -1556 106 -1552
rect 142 -1553 146 -1549
rect 436 -1550 440 -1546
rect 436 -1558 440 -1554
rect 285 -1564 289 -1560
rect 234 -1576 238 -1572
rect 436 -1566 440 -1562
rect 436 -1574 440 -1570
rect 437 -1638 441 -1634
rect 13 -1659 17 -1655
rect 50 -1659 54 -1655
rect 83 -1656 87 -1652
rect 437 -1646 441 -1642
rect 437 -1654 441 -1650
rect 102 -1674 106 -1670
rect 102 -1686 106 -1682
rect 224 -1669 228 -1665
rect 341 -1669 345 -1665
rect 224 -1677 228 -1673
rect 437 -1662 441 -1658
rect 437 -1670 441 -1666
rect 102 -1697 106 -1693
rect 142 -1694 146 -1690
rect 433 -1741 437 -1737
rect 433 -1749 437 -1745
rect 433 -1757 437 -1753
rect 433 -1765 437 -1761
rect 433 -1773 437 -1769
rect 433 -1781 437 -1777
rect 430 -1834 434 -1830
rect 430 -1842 434 -1838
rect 430 -1850 434 -1846
rect 430 -1858 434 -1854
rect 430 -1866 434 -1862
rect 430 -1874 434 -1870
rect 13 -1988 17 -1984
rect 50 -1988 54 -1984
rect 83 -1985 87 -1981
rect 102 -2003 106 -1999
rect 102 -2015 106 -2011
rect 102 -2026 106 -2022
rect 142 -2023 146 -2019
<< metal1 >>
rect 265 100 308 101
rect 269 96 308 100
rect 9 90 155 94
rect 9 62 12 90
rect 17 74 21 77
rect 39 62 42 90
rect 50 82 61 87
rect 54 74 59 82
rect 58 70 59 74
rect 79 62 82 90
rect 105 82 109 90
rect 87 77 91 80
rect 94 66 100 69
rect 97 59 100 66
rect 97 55 106 59
rect 28 43 32 46
rect 58 42 62 46
rect 101 43 106 47
rect 101 42 105 43
rect 58 38 105 42
rect 28 33 32 38
rect 58 33 62 38
rect 101 36 105 38
rect 121 39 125 62
rect 145 66 149 90
rect 260 87 285 92
rect 225 83 264 87
rect 153 39 157 46
rect 101 32 106 36
rect 121 35 146 39
rect 153 35 163 39
rect 121 29 125 35
rect 153 32 157 35
rect 12 5 16 23
rect 42 5 47 23
rect 105 5 109 19
rect 145 5 149 22
rect 225 19 229 83
rect 268 57 272 63
rect 283 57 287 63
rect 268 53 287 57
rect 268 50 272 53
rect 236 46 240 50
rect 244 19 248 26
rect 275 46 279 53
rect 283 44 287 53
rect 260 19 264 40
rect 291 57 295 63
rect 303 57 308 96
rect 291 53 308 57
rect 291 44 295 53
rect 483 49 487 58
rect 434 42 436 46
rect 448 45 457 49
rect 483 45 490 49
rect 434 34 436 38
rect 448 33 452 45
rect 483 41 487 45
rect 477 37 487 41
rect 452 29 457 33
rect 510 29 514 33
rect 288 19 292 27
rect 225 15 237 19
rect 244 15 292 19
rect 244 12 248 15
rect -4 0 0 5
rect 4 0 159 5
rect -4 -133 2 0
rect 236 -2 240 2
rect 7 -48 153 -44
rect 157 -48 161 -44
rect 7 -76 10 -48
rect 15 -64 19 -61
rect 37 -76 40 -48
rect 48 -56 59 -51
rect 52 -64 57 -56
rect 56 -68 57 -64
rect 77 -76 80 -48
rect 103 -56 107 -48
rect 92 -72 98 -69
rect 95 -79 98 -72
rect 95 -83 104 -79
rect 26 -95 30 -92
rect 56 -96 60 -92
rect 99 -95 104 -91
rect 99 -96 103 -95
rect 56 -100 103 -96
rect 26 -105 30 -100
rect 56 -105 60 -100
rect 99 -102 103 -100
rect 119 -99 123 -76
rect 143 -72 147 -48
rect 483 -48 487 -39
rect 338 -53 342 -49
rect 274 -71 278 -62
rect 225 -78 227 -74
rect 239 -75 248 -71
rect 274 -75 281 -71
rect 434 -55 436 -51
rect 448 -52 457 -48
rect 483 -52 490 -48
rect 434 -63 436 -59
rect 448 -64 452 -52
rect 483 -56 487 -52
rect 477 -60 487 -56
rect 452 -68 457 -64
rect 510 -68 514 -64
rect 225 -86 227 -82
rect 239 -87 243 -75
rect 274 -79 278 -75
rect 268 -83 278 -79
rect 346 -80 350 -73
rect 331 -84 339 -80
rect 346 -84 360 -80
rect 346 -87 350 -84
rect 243 -91 248 -87
rect 301 -91 305 -87
rect 151 -99 155 -92
rect 99 -106 104 -102
rect 119 -103 144 -99
rect 151 -103 162 -99
rect 338 -101 342 -97
rect 119 -109 123 -103
rect 151 -106 155 -103
rect 10 -133 14 -115
rect 40 -133 45 -115
rect 103 -133 107 -119
rect 143 -133 147 -116
rect -4 -138 -2 -133
rect 2 -138 157 -133
rect -4 -274 2 -138
rect 265 -183 308 -182
rect 7 -189 153 -185
rect 157 -189 161 -185
rect 269 -187 308 -183
rect 7 -217 10 -189
rect 15 -205 19 -202
rect 37 -217 40 -189
rect 48 -197 59 -192
rect 52 -205 57 -197
rect 56 -209 57 -205
rect 77 -217 80 -189
rect 103 -197 107 -189
rect 92 -213 98 -210
rect 95 -220 98 -213
rect 95 -224 104 -220
rect 26 -236 30 -233
rect 56 -237 60 -233
rect 99 -236 104 -232
rect 99 -237 103 -236
rect 56 -241 103 -237
rect 26 -246 30 -241
rect 56 -246 60 -241
rect 99 -243 103 -241
rect 119 -240 123 -217
rect 143 -213 147 -189
rect 260 -196 285 -191
rect 225 -200 264 -196
rect 151 -240 155 -233
rect 99 -247 104 -243
rect 119 -244 144 -240
rect 151 -244 162 -240
rect 119 -250 123 -244
rect 151 -247 155 -244
rect 10 -274 14 -256
rect 40 -274 45 -256
rect 103 -274 107 -260
rect 143 -274 147 -257
rect 225 -264 229 -200
rect 268 -226 272 -220
rect 283 -226 287 -220
rect 268 -230 287 -226
rect 268 -233 272 -230
rect 236 -237 240 -233
rect 244 -264 248 -257
rect 275 -237 279 -230
rect 283 -239 287 -230
rect 260 -264 264 -243
rect 291 -226 295 -220
rect 303 -226 308 -187
rect 480 -212 484 -203
rect 431 -219 433 -215
rect 445 -216 454 -212
rect 480 -216 487 -212
rect 291 -230 308 -226
rect 431 -227 433 -223
rect 445 -228 449 -216
rect 480 -220 484 -216
rect 474 -224 484 -220
rect 291 -239 295 -230
rect 449 -232 454 -228
rect 507 -232 511 -228
rect 288 -264 292 -256
rect 225 -268 237 -264
rect 244 -268 292 -264
rect 244 -271 248 -268
rect -4 -279 -2 -274
rect 2 -279 157 -274
rect -4 -416 2 -279
rect 474 -278 478 -269
rect 236 -285 240 -281
rect 425 -285 427 -281
rect 468 -282 481 -278
rect 425 -293 427 -289
rect 439 -290 448 -286
rect 425 -301 427 -297
rect 439 -302 443 -290
rect 474 -294 478 -282
rect 468 -298 478 -294
rect 443 -306 448 -302
rect 511 -306 516 -302
rect 7 -331 153 -327
rect 157 -331 161 -327
rect 7 -359 10 -331
rect 15 -347 19 -344
rect 37 -359 40 -331
rect 48 -339 59 -334
rect 52 -347 57 -339
rect 56 -351 57 -347
rect 77 -359 80 -331
rect 103 -339 107 -331
rect 92 -355 98 -352
rect 95 -362 98 -355
rect 95 -366 104 -362
rect 26 -378 30 -375
rect 56 -379 60 -375
rect 99 -378 104 -374
rect 99 -379 103 -378
rect 56 -383 103 -379
rect 26 -388 30 -383
rect 56 -388 60 -383
rect 99 -385 103 -383
rect 119 -382 123 -359
rect 143 -355 147 -331
rect 341 -341 345 -337
rect 274 -354 278 -345
rect 225 -361 227 -357
rect 239 -358 248 -354
rect 274 -358 281 -354
rect 225 -369 227 -365
rect 239 -370 243 -358
rect 274 -362 278 -358
rect 474 -353 478 -344
rect 425 -360 427 -356
rect 468 -357 481 -353
rect 268 -366 278 -362
rect 349 -368 353 -361
rect 425 -368 427 -364
rect 439 -365 448 -361
rect 243 -374 248 -370
rect 301 -374 305 -370
rect 334 -372 342 -368
rect 349 -372 363 -368
rect 349 -375 353 -372
rect 151 -382 155 -375
rect 99 -389 104 -385
rect 119 -386 144 -382
rect 151 -386 162 -382
rect 425 -376 427 -372
rect 439 -377 443 -365
rect 474 -369 478 -357
rect 468 -373 478 -369
rect 443 -381 448 -377
rect 511 -381 516 -377
rect 119 -392 123 -386
rect 151 -389 155 -386
rect 10 -416 14 -398
rect 40 -416 45 -398
rect 341 -389 345 -385
rect 103 -416 107 -402
rect 143 -416 147 -399
rect -4 -421 -2 -416
rect 2 -421 157 -416
rect -4 -603 2 -421
rect 488 -486 492 -477
rect 439 -493 441 -489
rect 453 -490 462 -486
rect 488 -490 495 -486
rect 439 -501 441 -497
rect 453 -502 457 -490
rect 488 -494 492 -490
rect 482 -498 492 -494
rect 457 -506 462 -502
rect 515 -506 519 -502
rect 265 -512 308 -511
rect 7 -518 153 -514
rect 157 -518 161 -514
rect 269 -516 308 -512
rect 7 -546 10 -518
rect 15 -534 19 -531
rect 37 -546 40 -518
rect 48 -526 59 -521
rect 52 -534 57 -526
rect 56 -538 57 -534
rect 77 -546 80 -518
rect 103 -526 107 -518
rect 92 -542 98 -539
rect 95 -549 98 -542
rect 95 -553 104 -549
rect 26 -565 30 -562
rect 56 -566 60 -562
rect 99 -565 104 -561
rect 99 -566 103 -565
rect 56 -570 103 -566
rect 26 -575 30 -570
rect 56 -575 60 -570
rect 99 -572 103 -570
rect 119 -569 123 -546
rect 143 -542 147 -518
rect 260 -525 285 -520
rect 225 -529 264 -525
rect 151 -569 155 -562
rect 99 -576 104 -572
rect 119 -573 144 -569
rect 151 -573 162 -569
rect 119 -579 123 -573
rect 151 -576 155 -573
rect 10 -603 14 -585
rect 40 -603 45 -585
rect 103 -603 107 -589
rect 143 -603 147 -586
rect 225 -593 229 -529
rect 268 -555 272 -549
rect 283 -555 287 -549
rect 268 -559 287 -555
rect 268 -562 272 -559
rect 236 -566 240 -562
rect 244 -593 248 -586
rect 275 -566 279 -559
rect 283 -568 287 -559
rect 260 -593 264 -572
rect 291 -555 295 -549
rect 303 -555 308 -516
rect 482 -552 486 -543
rect 291 -559 308 -555
rect 433 -559 435 -555
rect 476 -556 489 -552
rect 291 -568 295 -559
rect 433 -567 435 -563
rect 447 -564 456 -560
rect 433 -575 435 -571
rect 447 -576 451 -564
rect 482 -568 486 -556
rect 476 -572 486 -568
rect 451 -580 456 -576
rect 519 -580 524 -576
rect 288 -593 292 -585
rect 225 -597 237 -593
rect 244 -597 292 -593
rect 244 -600 248 -597
rect -4 -608 -2 -603
rect 2 -608 157 -603
rect -4 -745 2 -608
rect 236 -614 240 -610
rect 482 -634 486 -624
rect 433 -641 435 -637
rect 447 -638 456 -634
rect 482 -638 489 -634
rect 433 -649 435 -645
rect 447 -650 451 -638
rect 482 -642 486 -638
rect 476 -646 486 -642
rect 7 -660 153 -656
rect 157 -660 161 -656
rect 433 -657 435 -653
rect 447 -654 456 -650
rect 7 -688 10 -660
rect 15 -676 19 -673
rect 37 -688 40 -660
rect 48 -668 59 -663
rect 52 -676 57 -668
rect 56 -680 57 -676
rect 77 -688 80 -660
rect 103 -668 107 -660
rect 92 -684 98 -681
rect 95 -691 98 -684
rect 95 -695 104 -691
rect 26 -707 30 -704
rect 56 -708 60 -704
rect 99 -707 104 -703
rect 99 -708 103 -707
rect 56 -712 103 -708
rect 26 -717 30 -712
rect 56 -717 60 -712
rect 99 -714 103 -712
rect 119 -711 123 -688
rect 143 -684 147 -660
rect 341 -667 345 -663
rect 433 -665 435 -661
rect 447 -666 451 -654
rect 482 -658 486 -646
rect 476 -662 486 -658
rect 274 -683 278 -674
rect 225 -690 227 -686
rect 239 -687 248 -683
rect 274 -687 281 -683
rect 451 -670 456 -666
rect 529 -670 534 -666
rect 225 -698 227 -694
rect 239 -699 243 -687
rect 274 -691 278 -687
rect 268 -695 278 -691
rect 349 -694 353 -687
rect 334 -698 342 -694
rect 349 -698 363 -694
rect 243 -703 248 -699
rect 301 -703 305 -699
rect 349 -701 353 -698
rect 151 -711 155 -704
rect 99 -718 104 -714
rect 119 -715 144 -711
rect 151 -715 162 -711
rect 341 -715 345 -711
rect 119 -721 123 -715
rect 151 -718 155 -715
rect 10 -745 14 -727
rect 40 -745 45 -727
rect 483 -724 487 -714
rect 103 -745 107 -731
rect 143 -745 147 -728
rect 434 -731 436 -727
rect 448 -728 457 -724
rect 483 -728 490 -724
rect 434 -739 436 -735
rect 448 -740 452 -728
rect 483 -732 487 -728
rect 477 -736 487 -732
rect -4 -750 -2 -745
rect 2 -750 157 -745
rect 434 -747 436 -743
rect 448 -744 457 -740
rect -4 -1093 2 -750
rect 434 -755 436 -751
rect 448 -756 452 -744
rect 483 -748 487 -736
rect 477 -752 487 -748
rect 452 -760 457 -756
rect 530 -760 535 -756
rect 490 -900 494 -891
rect 441 -907 443 -903
rect 455 -904 464 -900
rect 490 -904 497 -900
rect 441 -915 443 -911
rect 455 -916 459 -904
rect 490 -908 494 -904
rect 484 -912 494 -908
rect 459 -920 464 -916
rect 517 -920 521 -916
rect 484 -966 488 -957
rect 435 -973 437 -969
rect 478 -970 491 -966
rect 435 -981 437 -977
rect 449 -978 458 -974
rect 435 -989 437 -985
rect 449 -990 453 -978
rect 484 -982 488 -970
rect 478 -986 488 -982
rect 453 -994 458 -990
rect 521 -994 526 -990
rect 263 -1001 306 -1000
rect 7 -1008 153 -1004
rect 157 -1008 161 -1004
rect 267 -1005 306 -1001
rect 7 -1036 10 -1008
rect 15 -1024 19 -1021
rect 37 -1036 40 -1008
rect 48 -1016 59 -1011
rect 52 -1024 57 -1016
rect 56 -1028 57 -1024
rect 77 -1036 80 -1008
rect 103 -1016 107 -1008
rect 92 -1032 98 -1029
rect 95 -1039 98 -1032
rect 95 -1043 104 -1039
rect 26 -1055 30 -1052
rect 56 -1056 60 -1052
rect 99 -1055 104 -1051
rect 99 -1056 103 -1055
rect 56 -1060 103 -1056
rect 26 -1065 30 -1060
rect 56 -1065 60 -1060
rect 99 -1062 103 -1060
rect 119 -1059 123 -1036
rect 143 -1032 147 -1008
rect 258 -1014 283 -1009
rect 223 -1018 262 -1014
rect 151 -1059 155 -1052
rect 99 -1066 104 -1062
rect 119 -1063 144 -1059
rect 151 -1063 162 -1059
rect 119 -1069 123 -1063
rect 151 -1066 155 -1063
rect 10 -1093 14 -1075
rect 40 -1093 45 -1075
rect 103 -1093 107 -1079
rect 143 -1093 147 -1076
rect 223 -1082 227 -1018
rect 266 -1044 270 -1038
rect 281 -1044 285 -1038
rect 266 -1048 285 -1044
rect 266 -1051 270 -1048
rect 234 -1055 238 -1051
rect 242 -1082 246 -1075
rect 273 -1055 277 -1048
rect 281 -1057 285 -1048
rect 258 -1082 262 -1061
rect 289 -1044 293 -1038
rect 301 -1044 306 -1005
rect 289 -1048 306 -1044
rect 484 -1048 488 -1038
rect 289 -1057 293 -1048
rect 435 -1055 437 -1051
rect 449 -1052 458 -1048
rect 484 -1052 491 -1048
rect 435 -1063 437 -1059
rect 449 -1064 453 -1052
rect 484 -1056 488 -1052
rect 478 -1060 488 -1056
rect 435 -1071 437 -1067
rect 449 -1068 458 -1064
rect 286 -1082 290 -1074
rect 435 -1079 437 -1075
rect 223 -1086 235 -1082
rect 242 -1086 290 -1082
rect 449 -1080 453 -1068
rect 484 -1072 488 -1060
rect 478 -1076 488 -1072
rect 453 -1084 458 -1080
rect 531 -1084 536 -1080
rect 242 -1089 246 -1086
rect -4 -1098 -2 -1093
rect 2 -1098 157 -1093
rect -4 -1234 2 -1098
rect 234 -1103 238 -1099
rect 485 -1135 489 -1126
rect 479 -1139 492 -1135
rect 436 -1143 438 -1139
rect 5 -1149 151 -1145
rect 155 -1149 159 -1145
rect 452 -1147 465 -1143
rect 5 -1177 8 -1149
rect 13 -1165 17 -1162
rect 35 -1177 38 -1149
rect 46 -1157 57 -1152
rect 50 -1165 55 -1157
rect 54 -1169 55 -1165
rect 75 -1177 78 -1149
rect 101 -1157 105 -1149
rect 90 -1173 96 -1170
rect 93 -1180 96 -1173
rect 93 -1184 102 -1180
rect 24 -1196 28 -1193
rect 54 -1197 58 -1193
rect 97 -1196 102 -1192
rect 97 -1197 101 -1196
rect 54 -1201 101 -1197
rect 24 -1206 28 -1201
rect 54 -1206 58 -1201
rect 97 -1203 101 -1201
rect 117 -1200 121 -1177
rect 141 -1173 145 -1149
rect 340 -1152 344 -1148
rect 436 -1151 438 -1147
rect 272 -1172 276 -1163
rect 436 -1159 438 -1155
rect 452 -1159 456 -1147
rect 485 -1151 489 -1139
rect 479 -1155 489 -1151
rect 452 -1163 465 -1159
rect 436 -1167 438 -1163
rect 223 -1179 225 -1175
rect 237 -1176 246 -1172
rect 272 -1176 279 -1172
rect 223 -1187 225 -1183
rect 237 -1188 241 -1176
rect 272 -1180 276 -1176
rect 348 -1179 352 -1172
rect 436 -1175 438 -1171
rect 452 -1175 456 -1163
rect 485 -1167 489 -1155
rect 479 -1171 489 -1167
rect 456 -1179 465 -1175
rect 542 -1179 549 -1175
rect 266 -1184 276 -1180
rect 333 -1183 341 -1179
rect 348 -1183 362 -1179
rect 348 -1186 352 -1183
rect 241 -1192 246 -1188
rect 299 -1192 303 -1188
rect 149 -1200 153 -1193
rect 340 -1200 344 -1196
rect 97 -1207 102 -1203
rect 117 -1204 142 -1200
rect 149 -1204 160 -1200
rect 117 -1210 121 -1204
rect 149 -1207 153 -1204
rect 8 -1234 12 -1216
rect 38 -1234 43 -1216
rect 101 -1234 105 -1220
rect 141 -1234 145 -1217
rect 484 -1219 488 -1210
rect 478 -1223 491 -1219
rect 435 -1227 437 -1223
rect 451 -1231 464 -1227
rect 0 -1239 155 -1234
rect 435 -1235 437 -1231
rect -4 -1378 2 -1239
rect 435 -1243 437 -1239
rect 451 -1243 455 -1231
rect 484 -1235 488 -1223
rect 478 -1239 488 -1235
rect 451 -1247 464 -1243
rect 435 -1251 437 -1247
rect 435 -1259 437 -1255
rect 451 -1259 455 -1247
rect 484 -1251 488 -1239
rect 478 -1255 488 -1251
rect 455 -1263 464 -1259
rect 541 -1263 548 -1259
rect -9 -1382 2 -1378
rect -4 -1583 2 -1382
rect 489 -1395 493 -1386
rect 440 -1402 442 -1398
rect 454 -1399 463 -1395
rect 489 -1399 496 -1395
rect 440 -1410 442 -1406
rect 454 -1411 458 -1399
rect 489 -1403 493 -1399
rect 483 -1407 493 -1403
rect 458 -1415 463 -1411
rect 516 -1415 520 -1411
rect 483 -1461 487 -1452
rect 434 -1468 436 -1464
rect 477 -1465 490 -1461
rect 434 -1476 436 -1472
rect 448 -1473 457 -1469
rect 434 -1484 436 -1480
rect 448 -1485 452 -1473
rect 483 -1477 487 -1465
rect 477 -1481 487 -1477
rect 452 -1489 457 -1485
rect 520 -1489 525 -1485
rect 262 -1491 305 -1490
rect 5 -1498 151 -1494
rect 155 -1498 159 -1494
rect 266 -1495 305 -1491
rect 5 -1526 8 -1498
rect 13 -1514 17 -1511
rect 35 -1526 38 -1498
rect 46 -1506 57 -1501
rect 50 -1514 55 -1506
rect 54 -1518 55 -1514
rect 75 -1526 78 -1498
rect 101 -1506 105 -1498
rect 83 -1511 88 -1506
rect 90 -1522 96 -1519
rect 93 -1529 96 -1522
rect 93 -1533 102 -1529
rect 24 -1545 28 -1542
rect 54 -1546 58 -1542
rect 97 -1545 102 -1541
rect 97 -1546 101 -1545
rect 54 -1550 101 -1546
rect 24 -1555 28 -1550
rect 54 -1555 58 -1550
rect 97 -1552 101 -1550
rect 117 -1549 121 -1526
rect 141 -1522 145 -1498
rect 257 -1504 282 -1499
rect 222 -1508 261 -1504
rect 149 -1549 153 -1542
rect 97 -1556 102 -1552
rect 117 -1553 142 -1549
rect 149 -1553 160 -1549
rect 117 -1559 121 -1553
rect 149 -1556 153 -1553
rect 8 -1583 12 -1565
rect 38 -1583 43 -1565
rect 101 -1583 105 -1569
rect 141 -1583 145 -1566
rect 222 -1572 226 -1508
rect 265 -1534 269 -1528
rect 280 -1534 284 -1528
rect 265 -1538 284 -1534
rect 265 -1541 269 -1538
rect 233 -1545 237 -1541
rect 241 -1572 245 -1565
rect 272 -1545 276 -1538
rect 280 -1547 284 -1538
rect 257 -1572 261 -1551
rect 288 -1534 292 -1528
rect 300 -1534 305 -1495
rect 288 -1538 305 -1534
rect 288 -1547 292 -1538
rect 483 -1543 487 -1533
rect 434 -1550 436 -1546
rect 448 -1547 457 -1543
rect 483 -1547 490 -1543
rect 434 -1558 436 -1554
rect 448 -1559 452 -1547
rect 483 -1551 487 -1547
rect 477 -1555 487 -1551
rect 285 -1572 289 -1564
rect 434 -1566 436 -1562
rect 448 -1563 457 -1559
rect 222 -1576 234 -1572
rect 241 -1576 289 -1572
rect 434 -1574 436 -1570
rect 448 -1575 452 -1563
rect 483 -1567 487 -1555
rect 477 -1571 487 -1567
rect 241 -1579 245 -1576
rect 452 -1579 457 -1575
rect 530 -1579 535 -1575
rect 0 -1588 155 -1583
rect -4 -1724 2 -1588
rect 233 -1593 237 -1589
rect 484 -1630 488 -1621
rect 478 -1634 491 -1630
rect 5 -1639 151 -1635
rect 155 -1639 159 -1635
rect 340 -1638 344 -1634
rect 435 -1638 437 -1634
rect 5 -1667 8 -1639
rect 13 -1655 17 -1652
rect 35 -1667 38 -1639
rect 46 -1647 57 -1642
rect 50 -1655 55 -1647
rect 54 -1659 55 -1655
rect 75 -1667 78 -1639
rect 101 -1647 105 -1639
rect 90 -1663 96 -1660
rect 93 -1670 96 -1663
rect 93 -1674 102 -1670
rect 24 -1686 28 -1683
rect 54 -1687 58 -1683
rect 97 -1686 102 -1682
rect 97 -1687 101 -1686
rect 54 -1691 101 -1687
rect 24 -1696 28 -1691
rect 54 -1696 58 -1691
rect 97 -1693 101 -1691
rect 117 -1690 121 -1667
rect 141 -1663 145 -1639
rect 271 -1662 275 -1653
rect 451 -1642 464 -1638
rect 435 -1646 437 -1642
rect 435 -1654 437 -1650
rect 451 -1654 455 -1642
rect 484 -1646 488 -1634
rect 478 -1650 488 -1646
rect 451 -1658 464 -1654
rect 222 -1669 224 -1665
rect 236 -1666 245 -1662
rect 271 -1666 278 -1662
rect 348 -1665 352 -1658
rect 435 -1662 437 -1658
rect 222 -1677 224 -1673
rect 236 -1678 240 -1666
rect 271 -1670 275 -1666
rect 333 -1669 341 -1665
rect 348 -1669 362 -1665
rect 265 -1674 275 -1670
rect 348 -1672 352 -1669
rect 435 -1670 437 -1666
rect 451 -1670 455 -1658
rect 484 -1662 488 -1650
rect 478 -1666 488 -1662
rect 240 -1682 245 -1678
rect 298 -1682 302 -1678
rect 455 -1674 464 -1670
rect 541 -1674 548 -1670
rect 149 -1690 153 -1683
rect 340 -1686 344 -1682
rect 97 -1697 102 -1693
rect 117 -1694 142 -1690
rect 149 -1694 160 -1690
rect 117 -1700 121 -1694
rect 149 -1697 153 -1694
rect 8 -1724 12 -1706
rect 38 -1724 43 -1706
rect 101 -1724 105 -1710
rect 141 -1724 145 -1707
rect 0 -1729 155 -1724
rect -4 -2053 2 -1729
rect 480 -1734 484 -1724
rect 431 -1741 433 -1737
rect 445 -1738 454 -1734
rect 480 -1738 487 -1734
rect 431 -1749 433 -1745
rect 445 -1750 449 -1738
rect 480 -1742 484 -1738
rect 474 -1746 484 -1742
rect 431 -1757 433 -1753
rect 445 -1754 454 -1750
rect 431 -1765 433 -1761
rect 445 -1766 449 -1754
rect 480 -1758 484 -1746
rect 474 -1762 484 -1758
rect 431 -1773 433 -1769
rect 445 -1770 454 -1766
rect 431 -1781 433 -1777
rect 445 -1782 449 -1770
rect 480 -1774 484 -1762
rect 474 -1778 484 -1774
rect 449 -1786 454 -1782
rect 547 -1786 552 -1782
rect 477 -1827 481 -1817
rect 428 -1834 430 -1830
rect 442 -1831 451 -1827
rect 477 -1831 484 -1827
rect 428 -1842 430 -1838
rect 442 -1843 446 -1831
rect 477 -1835 481 -1831
rect 471 -1839 481 -1835
rect 428 -1850 430 -1846
rect 442 -1847 451 -1843
rect 428 -1858 430 -1854
rect 442 -1859 446 -1847
rect 477 -1851 481 -1839
rect 471 -1855 481 -1851
rect 428 -1866 430 -1862
rect 442 -1863 451 -1859
rect 428 -1874 430 -1870
rect 442 -1875 446 -1863
rect 477 -1867 481 -1855
rect 471 -1871 481 -1867
rect 446 -1879 451 -1875
rect 544 -1879 549 -1875
rect 5 -1968 151 -1964
rect 155 -1968 159 -1964
rect 5 -1996 8 -1968
rect 13 -1984 17 -1981
rect 35 -1996 38 -1968
rect 46 -1976 57 -1971
rect 50 -1984 55 -1976
rect 54 -1988 55 -1984
rect 75 -1996 78 -1968
rect 101 -1976 105 -1968
rect 90 -1992 96 -1989
rect 93 -1999 96 -1992
rect 93 -2003 102 -1999
rect 24 -2015 28 -2012
rect 54 -2016 58 -2012
rect 97 -2015 102 -2011
rect 97 -2016 101 -2015
rect 54 -2020 101 -2016
rect 24 -2025 28 -2020
rect 54 -2025 58 -2020
rect 97 -2022 101 -2020
rect 117 -2019 121 -1996
rect 141 -1992 145 -1968
rect 149 -2019 153 -2012
rect 97 -2026 102 -2022
rect 117 -2023 142 -2019
rect 149 -2023 160 -2019
rect 117 -2029 121 -2023
rect 149 -2026 153 -2023
rect 8 -2053 12 -2035
rect 38 -2053 43 -2035
rect 101 -2053 105 -2039
rect 141 -2053 145 -2036
rect 0 -2058 155 -2053
<< pm12contact >>
rect 25 70 30 75
rect 45 70 50 75
rect 117 10 122 15
rect 23 -68 28 -63
rect 43 -68 48 -63
rect 115 -128 120 -123
rect 23 -209 28 -204
rect 43 -209 48 -204
rect 115 -269 120 -264
rect 23 -351 28 -346
rect 43 -351 48 -346
rect 115 -411 120 -406
rect 23 -538 28 -533
rect 43 -538 48 -533
rect 115 -598 120 -593
rect 23 -680 28 -675
rect 43 -680 48 -675
rect 115 -740 120 -735
rect 23 -1028 28 -1023
rect 43 -1028 48 -1023
rect 115 -1088 120 -1083
rect 21 -1169 26 -1164
rect 41 -1169 46 -1164
rect 113 -1229 118 -1224
rect 21 -1518 26 -1513
rect 41 -1518 46 -1513
rect 113 -1578 118 -1573
rect 21 -1659 26 -1654
rect 41 -1659 46 -1654
rect 113 -1719 118 -1714
rect 21 -1988 26 -1983
rect 41 -1988 46 -1983
rect 113 -2048 118 -2043
<< metal2 >>
rect 0 80 28 83
rect 0 48 3 80
rect 24 77 28 80
rect 24 75 50 77
rect 24 74 25 75
rect 30 74 45 75
rect -28 42 3 48
rect -28 -78 -22 42
rect 0 12 3 42
rect 0 10 117 12
rect 0 9 121 10
rect -2 -58 26 -55
rect -2 -78 1 -58
rect 22 -61 26 -58
rect 22 -63 48 -61
rect 22 -64 23 -63
rect 28 -64 43 -63
rect -28 -84 1 -78
rect -28 -244 -22 -84
rect -2 -126 1 -84
rect -2 -128 115 -126
rect -2 -129 119 -128
rect -2 -199 26 -196
rect -2 -244 1 -199
rect 22 -202 26 -199
rect 22 -204 48 -202
rect 22 -205 23 -204
rect 28 -205 43 -204
rect -28 -250 1 -244
rect -28 -373 -22 -250
rect -2 -267 1 -250
rect -2 -269 115 -267
rect -2 -270 119 -269
rect -2 -341 26 -338
rect -2 -373 1 -341
rect 22 -344 26 -341
rect 22 -346 48 -344
rect 22 -347 23 -346
rect 28 -347 43 -346
rect -28 -379 1 -373
rect -28 -565 -22 -379
rect -2 -409 1 -379
rect -2 -411 115 -409
rect -2 -412 119 -411
rect -2 -528 26 -525
rect -2 -565 1 -528
rect 22 -531 26 -528
rect 22 -533 48 -531
rect 22 -534 23 -533
rect 28 -534 43 -533
rect -28 -571 1 -565
rect -28 -699 -22 -571
rect -2 -596 1 -571
rect -2 -598 115 -596
rect -2 -599 119 -598
rect -2 -670 26 -667
rect -2 -699 1 -670
rect 22 -673 26 -670
rect 22 -675 48 -673
rect 22 -676 23 -675
rect 28 -676 43 -675
rect -28 -705 1 -699
rect -28 -931 -22 -705
rect -2 -738 1 -705
rect -2 -740 115 -738
rect -2 -741 119 -740
rect -42 -936 -22 -931
rect -28 -1045 -22 -936
rect -2 -1018 26 -1015
rect -2 -1045 1 -1018
rect 22 -1021 26 -1018
rect 22 -1023 48 -1021
rect 22 -1024 23 -1023
rect 28 -1024 43 -1023
rect -28 -1051 1 -1045
rect -28 -1199 -22 -1051
rect -2 -1086 1 -1051
rect -2 -1088 115 -1086
rect -2 -1089 119 -1088
rect -4 -1159 24 -1156
rect -4 -1199 -1 -1159
rect 20 -1162 24 -1159
rect 20 -1164 46 -1162
rect 20 -1165 21 -1164
rect 26 -1165 41 -1164
rect -28 -1205 0 -1199
rect -28 -1555 -22 -1205
rect -4 -1227 -1 -1205
rect -4 -1229 113 -1227
rect -4 -1230 117 -1229
rect -4 -1508 24 -1505
rect -4 -1555 -1 -1508
rect 20 -1511 24 -1508
rect 20 -1513 46 -1511
rect 20 -1514 21 -1513
rect 26 -1514 41 -1513
rect -28 -1561 0 -1555
rect -28 -1686 -22 -1561
rect -4 -1576 -1 -1561
rect -4 -1578 113 -1576
rect -4 -1579 117 -1578
rect -4 -1649 24 -1646
rect -4 -1686 -1 -1649
rect 20 -1652 24 -1649
rect 20 -1654 46 -1652
rect 20 -1655 21 -1654
rect 26 -1655 41 -1654
rect -28 -1692 0 -1686
rect -28 -2009 -22 -1692
rect -4 -1717 -1 -1692
rect -4 -1719 113 -1717
rect -4 -1720 117 -1719
rect -4 -1978 24 -1975
rect -4 -2009 -1 -1978
rect 20 -1981 24 -1978
rect 20 -1983 46 -1981
rect 20 -1984 21 -1983
rect 26 -1984 41 -1983
rect -28 -2015 0 -2009
rect -4 -2046 -1 -2015
rect -4 -2048 113 -2046
rect -4 -2049 117 -2048
<< m3contact >>
rect 83 -1511 88 -1506
<< m123contact >>
rect 45 82 50 87
rect 87 80 92 85
rect 28 38 33 43
rect 43 -56 48 -51
rect 85 -61 90 -56
rect 26 -100 31 -95
rect 43 -197 48 -192
rect 85 -202 90 -197
rect 26 -241 31 -236
rect 43 -339 48 -334
rect 85 -344 90 -339
rect 26 -383 31 -378
rect 43 -526 48 -521
rect 85 -531 90 -526
rect 26 -570 31 -565
rect 43 -668 48 -663
rect 85 -673 90 -668
rect 26 -712 31 -707
rect 43 -1016 48 -1011
rect 85 -1021 90 -1016
rect 26 -1060 31 -1055
rect 41 -1157 46 -1152
rect 83 -1162 88 -1157
rect 24 -1201 29 -1196
rect 41 -1506 46 -1501
rect 24 -1550 29 -1545
rect 41 -1647 46 -1642
rect 83 -1652 88 -1647
rect 24 -1691 29 -1686
rect 41 -1976 46 -1971
rect 83 -1981 88 -1976
rect 24 -2020 29 -2015
<< metal3 >>
rect 159 90 190 94
rect 35 82 45 87
rect 35 43 38 82
rect 75 80 87 83
rect 33 38 39 43
rect 33 -56 43 -51
rect 33 -95 36 -56
rect 75 -58 78 80
rect 75 -61 85 -58
rect 31 -100 37 -95
rect 33 -197 43 -192
rect 33 -236 36 -197
rect 75 -199 78 -61
rect 75 -202 85 -199
rect 31 -241 37 -236
rect 33 -339 43 -334
rect 33 -378 36 -339
rect 75 -341 78 -202
rect 75 -344 85 -341
rect 31 -383 37 -378
rect 33 -526 43 -521
rect 33 -565 36 -526
rect 75 -528 78 -344
rect 75 -531 85 -528
rect 31 -570 37 -565
rect 33 -668 43 -663
rect 33 -707 36 -668
rect 75 -670 78 -531
rect 75 -673 85 -670
rect 31 -712 37 -707
rect 75 -881 78 -673
rect 63 -885 78 -881
rect 33 -1016 43 -1011
rect 33 -1055 36 -1016
rect 75 -1018 78 -885
rect 75 -1021 85 -1018
rect 31 -1060 37 -1055
rect 31 -1157 41 -1152
rect 31 -1196 34 -1157
rect 75 -1159 78 -1021
rect 75 -1162 83 -1159
rect 29 -1201 35 -1196
rect 31 -1506 41 -1501
rect 31 -1545 34 -1506
rect 75 -1508 78 -1162
rect 75 -1511 83 -1508
rect 29 -1550 35 -1545
rect 31 -1647 41 -1642
rect 31 -1686 34 -1647
rect 75 -1649 78 -1511
rect 75 -1652 83 -1649
rect 29 -1691 35 -1686
rect 31 -1976 41 -1971
rect 31 -2015 34 -1976
rect 75 -1978 78 -1652
rect 75 -1981 83 -1978
rect 29 -2020 35 -2015
rect 186 -2039 190 90
<< labels >>
rlabel metal1 17 74 21 77 1 a0
rlabel metal1 15 -64 19 -61 1 b0
rlabel metal1 15 -205 19 -202 1 a1
rlabel metal1 15 -347 19 -344 1 b1
rlabel metal1 15 -534 19 -531 1 a2
rlabel metal1 15 -676 19 -673 1 b2
rlabel metal1 15 -1024 19 -1021 1 a3
rlabel metal1 13 -1165 17 -1162 1 b3
rlabel metal1 13 -1514 17 -1511 1 a4
rlabel metal1 13 -1655 17 -1652 1 b4
rlabel metal1 13 -1984 17 -1981 1 c0
rlabel metal2 -42 -936 -28 -931 1 clk
rlabel metal3 63 -885 75 -881 1 rst
rlabel metal1 -9 -1382 -4 -1378 1 gnd
<< end >>
