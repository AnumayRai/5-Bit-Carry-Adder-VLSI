magic
tech scmos
timestamp 1763328877
<< nwell >>
rect 9 -46 49 -6
<< ntransistor >>
rect 56 -19 86 -17
rect 56 -27 86 -25
rect 56 -35 86 -33
<< ptransistor >>
rect 23 -19 43 -17
rect 23 -27 43 -25
rect 23 -35 43 -33
<< ndiffusion >>
rect 56 -17 86 -16
rect 56 -20 86 -19
rect 56 -25 86 -24
rect 56 -28 86 -27
rect 56 -33 86 -32
rect 56 -36 86 -35
<< pdiffusion >>
rect 23 -17 43 -16
rect 23 -20 43 -19
rect 23 -25 43 -24
rect 23 -28 43 -27
rect 23 -33 43 -32
rect 23 -36 43 -35
<< ndcontact >>
rect 56 -16 86 -12
rect 56 -24 86 -20
rect 56 -32 86 -28
rect 56 -40 86 -36
<< pdcontact >>
rect 23 -16 43 -12
rect 23 -24 43 -20
rect 23 -32 43 -28
rect 23 -40 43 -36
<< psubstratepcontact >>
rect 91 -40 95 -36
<< nsubstratencontact >>
rect 14 -40 18 -36
<< polysilicon >>
rect 6 -19 23 -17
rect 43 -19 56 -17
rect 86 -19 89 -17
rect 6 -27 23 -25
rect 43 -27 56 -25
rect 86 -27 89 -25
rect 6 -35 23 -33
rect 43 -35 56 -33
rect 86 -35 89 -33
<< polycontact >>
rect 2 -19 6 -15
rect 2 -27 6 -23
rect 2 -35 6 -31
<< metal1 >>
rect 49 -12 53 -3
rect 0 -19 2 -15
rect 43 -16 56 -12
rect 0 -27 2 -23
rect 14 -24 23 -20
rect 0 -35 2 -31
rect 14 -36 18 -24
rect 49 -28 53 -16
rect 43 -32 53 -28
rect 18 -40 23 -36
rect 86 -40 91 -36
<< labels >>
rlabel nsubstratencontact 14 -40 18 -36 7 vdd
rlabel metal1 0 -35 2 -33 3 a
rlabel metal1 0 -27 2 -25 3 b
rlabel metal1 0 -19 2 -17 3 c
rlabel metal1 49 -5 53 -3 5 vo
rlabel psubstratepcontact 91 -40 95 -36 7 gnd
<< end >>
