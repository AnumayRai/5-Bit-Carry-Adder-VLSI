magic
tech scmos
timestamp 1763239429
<< nwell >>
rect 0 0 24 37
<< ntransistor >>
rect 11 -18 13 -8
<< ptransistor >>
rect 11 6 13 26
<< ndiffusion >>
rect 10 -18 11 -8
rect 13 -18 14 -8
<< pdiffusion >>
rect 10 6 11 26
rect 13 6 14 26
<< ndcontact >>
rect 6 -18 10 -8
rect 14 -18 18 -8
<< pdcontact >>
rect 6 6 10 26
rect 14 6 18 26
<< psubstratepcontact >>
rect 6 -26 10 -22
<< nsubstratencontact >>
rect 6 30 10 34
<< polysilicon >>
rect 11 26 13 29
rect 11 -8 13 6
rect 11 -21 13 -18
<< polycontact >>
rect 7 -5 11 -1
<< metal1 >>
rect 6 26 10 30
rect 14 -1 18 6
rect -1 -5 7 -1
rect 14 -5 28 -1
rect 14 -8 18 -5
rect 6 -22 10 -18
<< labels >>
rlabel metal1 6 -23 10 -22 1 gnd
rlabel metal1 -1 -5 0 -1 3 a
rlabel metal1 26 -5 28 -1 7 b
rlabel metal1 6 31 10 33 5 vdd
<< end >>
