CLA with D Flip Flop
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

    
Vdd	vdd	gnd	'SUPPLY'
vclk clk gnd pulse 1.8 0 2ns 0ns 0ns 45ns 90ns
vrst rst gnd pulse 1.8 0 1ns 0ns 0ns 45ns 700ns


* A = 0 0 1 0 1  (a4..a0)
va0 a0 gnd 1.8
va1 a1 gnd 0
va2 a2 gnd 1.8
va3 a3 gnd 0
va4 a4 gnd 0

* B = 0 1 0 0 1  (b4..b0)
vb0 b0 gnd 1.8
vb1 b1 gnd 0
vb2 b2 gnd 0
vb3 b3 gnd 0
vb4 b4 gnd 0

* Cin
vc0 c0 gnd 0



.option scale=0.09u

M1000 q0 a_243_2# p0 Gnd cmosn w=10 l=2
+  ad=100 pd=60 as=100 ps=60
M1001 a_47_n92# clk vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=12674 ps=6230
M1002 a_17_n115# b0 gnd Gnd cmosn w=10 l=2
+  ad=130 pd=46 as=6700 ps=3470
M1003 a_17_n256# clk a_17_n233# vdd cmosp w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1004 q7 qb7 vdd vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1005 qb8 clk a_108_n1220# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=60 ps=32
M1006 a_110_n402# a_55_n398# gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1007 qb5 clk a_110_n119# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=60 ps=32
M1008 a_241_n1099# q8 vdd vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1009 a_279_n1185# q8 gnd Gnd cmosn w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1010 a_840_n663# p1 vdd vdd cmosp w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1011 a_873_n655# p0 a_873_n663# Gnd cmosn w=40 l=2
+  ad=240 pd=92 as=240 ps=92
M1012 qb0 a_57_23# vdd vdd cmosp w=20 l=2
+  ad=260 pd=66 as=0 ps=0
M1013 p0 q0 q5 vdd cmosp w=20 l=2
+  ad=200 pd=100 as=200 ps=100
M1014 q1 qb1 gnd Gnd cmosn w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1015 a_47_n375# clk vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1016 vdd p4 a_838_n1779# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=360 ps=156
M1017 qb6 a_55_n398# vdd vdd cmosp w=20 l=2
+  ad=260 pd=66 as=0 ps=0
M1018 qb3 clk a_110_n1079# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=60 ps=32
M1019 a_875_n1069# p1 a_875_n1077# Gnd cmosn w=40 l=2
+  ad=240 pd=92 as=240 ps=92
M1020 a_841_36# p0 a_874_36# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1021 a_55_n256# a_17_n256# a_47_n256# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=60 ps=32
M1022 a_848_n1667# p2 vdd vdd cmosp w=14 l=2
+  ad=238 pd=118 as=0 ps=0
M1023 q0 q5 p0 vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1024 vdd p1 a_840_n573# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1025 a_873_n573# g0 gnd Gnd cmosn w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1026 p3 q3 a_241_n1099# Gnd cmosn w=10 l=2
+  ad=100 pd=60 as=100 ps=60
M1027 g2 g2_bar vdd vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1028 a_849_n1172# qc0 vdd vdd cmosp w=14 l=2
+  ad=238 pd=118 as=0 ps=0
M1029 g4_bar q9 vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1030 a_281_n84# q5 gnd Gnd cmosn w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1031 a_17_n704# b2 vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1032 g2_bar q2 a_281_n696# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1033 a_110_n260# a_55_n256# gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1034 c2 a_838_n225# vdd vdd cmosp w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1035 a_1057_n246# g1_bar a_1057_n254# Gnd cmosn w=30 l=2
+  ad=180 pd=72 as=180 ps=72
M1036 a_842_n987# g1 vdd vdd cmosp w=20 l=2
+  ad=220 pd=102 as=0 ps=0
M1037 g4_bar q4 a_278_n1675# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1038 vdd a_847_n1408# cout vdd cmosp w=20 l=2
+  ad=0 pd=0 as=360 ps=156
M1039 a_55_n256# rst vdd vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1040 g1 g1_bar gnd Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1041 qc0 qbc0 gnd Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1042 qb4 a_53_n1565# vdd vdd cmosp w=20 l=2
+  ad=260 pd=66 as=0 ps=0
M1043 a_17_n115# clk a_17_n92# vdd cmosp w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1044 vdd p0 a_832_n299# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1045 a_17_n398# clk a_17_n375# vdd cmosp w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1046 a_281_n367# q6 gnd Gnd cmosn w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1047 c3 a_840_n573# vdd vdd cmosp w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1048 a_1066_n585# g2_bar a_1066_n593# Gnd cmosn w=40 l=2
+  ad=240 pd=92 as=240 ps=92
M1049 vdd p3 a_842_n1077# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=240 ps=104
M1050 vdd q1 g1_bar vdd cmosp w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1051 a_881_n913# g2 gnd Gnd cmosn w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1052 a_15_n2035# clk a_15_n2012# vdd cmosp w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1053 a_47_n727# clk gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1054 a_15_n1216# clk a_15_n1193# vdd cmosp w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1055 qb9 clk a_108_n1710# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=60 ps=32
M1056 a_875_n1659# p1 a_875_n1667# Gnd cmosn w=50 l=2
+  ad=300 pd=112 as=300 ps=112
M1057 a_1091_n1048# a_842_n1077# a_1091_n1056# Gnd cmosn w=50 l=2
+  ad=300 pd=112 as=300 ps=112
M1058 a_243_2# q5 vdd vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1059 q6 qb6 gnd Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1060 vdd p2 a_849_n1172# vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1061 a_871_n1771# p0 a_871_n1779# Gnd cmosn w=60 l=2
+  ad=360 pd=132 as=360 ps=132
M1062 a_865_n299# qc0 gnd Gnd cmosn w=30 l=2
+  ad=180 pd=72 as=0 ps=0
M1063 c1 a_841_36# a_970_n61# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1064 g0_bar q5 vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1065 a_55_n398# a_17_n398# a_47_n398# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=60 ps=32
M1066 p2 q2 a_243_n610# Gnd cmosn w=10 l=2
+  ad=100 pd=60 as=100 ps=60
M1067 q8 qb8 gnd Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1068 qb0 clk a_112_19# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=60 ps=32
M1069 a_840_n663# p2 a_873_n647# Gnd cmosn w=40 l=2
+  ad=200 pd=90 as=240 ps=92
M1070 a_45_n1542# clk vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1071 a_838_n1779# p1 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 a_1098_n1572# a_838_n1779# gnd Gnd cmosn w=60 l=2
+  ad=360 pd=132 as=0 ps=0
M1073 a_874_n1572# g1 gnd Gnd cmosn w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1074 a_19_23# a0 gnd Gnd cmosn w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1075 a_47_n562# clk vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1076 qb2 a_55_n585# vdd vdd cmosp w=20 l=2
+  ad=260 pd=66 as=0 ps=0
M1077 q3 qb3 gnd Gnd cmosn w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1078 a_55_n115# a_17_n115# a_47_n92# vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1079 c4 a_848_n913# vdd vdd cmosp w=14 l=2
+  ad=238 pd=118 as=0 ps=0
M1080 vdd p4 a_847_n1408# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1081 a_848_n1667# p4 a_875_n1643# Gnd cmosn w=50 l=2
+  ad=250 pd=110 as=300 ps=112
M1082 a_17_n1075# clk a_17_n1052# vdd cmosp w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1083 a_876_n1156# p1 a_876_n1164# Gnd cmosn w=50 l=2
+  ad=300 pd=112 as=300 ps=112
M1084 a_15_n1565# a4 gnd Gnd cmosn w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1085 q2 q7 p2 vdd cmosp w=20 l=2
+  ad=200 pd=100 as=200 ps=100
M1086 a_842_n987# p3 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 a_875_n979# p2 a_875_n987# Gnd cmosn w=30 l=2
+  ad=180 pd=72 as=180 ps=72
M1088 g3 g3_bar gnd Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1089 a_45_n2035# clk gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1090 a_871_n1747# p3 a_871_n1755# Gnd cmosn w=60 l=2
+  ad=360 pd=132 as=360 ps=132
M1091 a_838_n225# g0 vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1092 vdd a_841_36# c1 vdd cmosp w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1093 a_53_n2035# rst vdd vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1094 cout a_841_n1572# vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 a_841_n1572# p3 vdd vdd cmosp w=20 l=2
+  ad=240 pd=104 as=0 ps=0
M1096 c3 a_846_n499# a_1066_n577# Gnd cmosn w=40 l=2
+  ad=200 pd=90 as=240 ps=92
M1097 a_53_n1216# rst vdd vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1098 a_55_n256# a_17_n256# a_47_n233# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1099 a_842_n1077# g0 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 a_15_n1706# clk a_15_n1683# vdd cmosp w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1101 a_1098_n1548# g4_bar a_1098_n1556# Gnd cmosn w=60 l=2
+  ad=360 pd=132 as=360 ps=132
M1102 a_841_n1572# p4 a_874_n1556# Gnd cmosn w=40 l=2
+  ad=200 pd=90 as=240 ps=92
M1103 a_108_n1569# a_53_n1565# gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1104 a_47_n115# clk gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1105 a_17_n585# clk a_17_n562# vdd cmosp w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1106 vdd p3 a_841_n1482# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=220 ps=102
M1107 a_846_n499# p2 a_879_n499# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1108 a_110_n731# a_55_n727# gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1109 a_1091_n1032# a_842_n987# a_1091_n1040# Gnd cmosn w=50 l=2
+  ad=300 pd=112 as=300 ps=112
M1110 a_45_n1216# clk gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1111 a_841_n1482# p4 a_874_n1474# Gnd cmosn w=30 l=2
+  ad=150 pd=70 as=180 ps=72
M1112 q9 qb9 gnd Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1113 q2 qb2 gnd Gnd cmosn w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1114 a_55_n727# rst vdd vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1115 q3 a_241_n1099# p3 Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 qb7 a_55_n727# vdd vdd cmosp w=20 l=2
+  ad=260 pd=66 as=0 ps=0
M1117 a_19_46# a0 vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1118 q5 qb5 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 a_55_n585# a_17_n585# a_47_n585# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=60 ps=32
M1120 vdd p0 a_840_n663# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1121 a_873_n663# qc0 gnd Gnd cmosn w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 a_47_n1075# clk gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1123 p1 q1 q6 vdd cmosp w=20 l=2
+  ad=200 pd=100 as=200 ps=100
M1124 g2 g2_bar gnd Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1125 q4 qb4 vdd vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1126 a_47_n704# clk vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1127 a_55_n1075# rst vdd vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1128 a_53_n1565# a_15_n1565# a_45_n1565# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=60 ps=32
M1129 a_110_n589# a_55_n585# gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1130 a_840_n573# g0 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1131 vdd p1 a_848_n1667# vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 g4 g4_bar vdd vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1133 qb6 clk a_110_n402# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1134 vdd p3 a_848_n913# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1135 vdd a_842_n1077# c4 vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 a_55_n585# rst vdd vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1137 a_849_n1172# p3 a_876_n1148# Gnd cmosn w=50 l=2
+  ad=250 pd=110 as=300 ps=112
M1138 a_838_n225# p1 a_871_n225# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1139 a_55_n398# a_17_n398# a_47_n375# vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1140 a_281_n696# q7 gnd Gnd cmosn w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 q0 qb0 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1142 vdd g1_bar c2 vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1143 a_1057_n254# a_832_n299# gnd Gnd cmosn w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 qb8 a_53_n1216# vdd vdd cmosp w=20 l=2
+  ad=260 pd=66 as=0 ps=0
M1145 vdd a_225_n1179# g3_bar vdd cmosp w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1146 a_278_n1675# q9 gnd Gnd cmosn w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 a_53_n1706# rst vdd vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1148 a_240_n1589# q9 vdd vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1149 cout a_841_n1482# vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1150 a_49_23# clk gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1151 vdd g2_bar c3 vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1152 a_1066_n593# a_840_n663# gnd Gnd cmosn w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1153 a_842_n1077# p2 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1154 a_880_n1408# g3 gnd Gnd cmosn w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1155 cout a_847_n1408# a_1098_n1540# Gnd cmosn w=60 l=2
+  ad=300 pd=130 as=360 ps=132
M1156 a_17_n256# a1 gnd Gnd cmosn w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1157 g0 g0_bar vdd vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1158 a_842_n1077# p3 a_875_n1061# Gnd cmosn w=40 l=2
+  ad=200 pd=90 as=240 ps=92
M1159 a_45_n1706# clk gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1160 p4 q4 a_240_n1589# Gnd cmosn w=10 l=2
+  ad=100 pd=60 as=100 ps=60
M1161 qb1 clk a_110_n260# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1162 a_17_n727# clk a_17_n704# vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1163 a_848_n1667# p4 vdd vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 a_840_n573# p2 a_873_n565# Gnd cmosn w=30 l=2
+  ad=150 pd=70 as=180 ps=72
M1165 a_1091_n1056# a_849_n1172# gnd Gnd cmosn w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 a_15_n1542# a4 vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1167 a_849_n1172# p1 vdd vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 a_45_n2012# clk vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1169 a_871_n1779# qc0 gnd Gnd cmosn w=60 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 a_832_n299# qc0 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1171 a_45_n1193# clk vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1172 a_970_n61# g0_bar gnd Gnd cmosn w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 vdd p2 a_840_n663# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1174 q7 qb7 gnd Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1175 qb3 a_55_n1075# vdd vdd cmosp w=20 l=2
+  ad=260 pd=66 as=0 ps=0
M1176 a_55_n727# a_17_n727# a_47_n727# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1177 a_241_n1099# q8 gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1178 vdd p0 a_838_n1779# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 a_832_n299# p1 a_865_n291# Gnd cmosn w=30 l=2
+  ad=150 pd=70 as=180 ps=72
M1180 a_15_n2035# c0 gnd Gnd cmosn w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1181 a_243_n610# q7 gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1182 p3 q3 q8 vdd cmosp w=20 l=2
+  ad=200 pd=100 as=200 ps=100
M1183 vdd a_842_n987# c4 vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1184 a_875_n1643# p3 a_875_n1651# Gnd cmosn w=50 l=2
+  ad=0 pd=0 as=300 ps=112
M1185 qb9 a_53_n1706# vdd vdd cmosp w=20 l=2
+  ad=260 pd=66 as=0 ps=0
M1186 a_876_n1164# p0 a_876_n1172# Gnd cmosn w=50 l=2
+  ad=0 pd=0 as=300 ps=112
M1187 a_17_n398# b1 gnd Gnd cmosn w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1188 a_55_n585# a_17_n585# a_47_n562# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 vdd p2 a_842_n987# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1190 a_871_n1755# p2 a_871_n1763# Gnd cmosn w=60 l=2
+  ad=0 pd=0 as=360 ps=132
M1191 a_108_n2039# a_53_n2035# gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1192 c1 g0_bar vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1193 q1 qb1 vdd vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1194 a_47_n1052# clk vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1195 vdd a_848_n1667# cout vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1196 vdd p2 a_841_n1572# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 a_49_46# clk vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1198 q0 qb0 gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1199 g1_bar q1 a_281_n367# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1200 vdd a_846_n499# c3 vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1201 a_15_n1216# b3 gnd Gnd cmosn w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1202 a_838_n1779# p3 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1203 a_1098_n1556# a_841_n1572# a_1098_n1564# Gnd cmosn w=60 l=2
+  ad=0 pd=0 as=360 ps=132
M1204 a_874_n1556# p3 a_874_n1564# Gnd cmosn w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1205 a_53_n1565# a_15_n1565# a_45_n1542# vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1206 a_875_n1077# g0 gnd Gnd cmosn w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 vdd p2 a_846_n499# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1208 a_1091_n1040# g3_bar a_1091_n1048# Gnd cmosn w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 g4 g4_bar gnd Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1210 a_45_n1683# clk vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1211 a_841_n1482# g2 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 q3 q8 p3 vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1213 a_849_n1172# p3 vdd vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 a_874_n1474# p3 a_874_n1482# Gnd cmosn w=30 l=2
+  ad=0 pd=0 as=180 ps=72
M1215 q5 qb5 gnd Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1216 a_17_n1075# a3 gnd Gnd cmosn w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1217 a_108_n1220# a_53_n1216# gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1218 a_57_23# rst vdd vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1219 a_55_n115# a_17_n115# a_47_n115# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1220 g1 g1_bar vdd vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1221 p2 q2 q7 vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1222 qc0 qbc0 vdd vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1223 a_243_2# q5 gnd Gnd cmosn w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1224 a_840_n663# qc0 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1225 vdd q2 g2_bar vdd cmosp w=20 l=2
+  ad=0 pd=0 as=120 ps=52
M1226 a_53_n2035# a_15_n2035# a_45_n2035# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1227 a_17_n233# a1 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 qb7 clk a_110_n731# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1229 q8 qb8 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 a_879_n499# g1 gnd Gnd cmosn w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1231 a_110_n1079# a_55_n1075# gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 a_841_36# qc0 vdd vdd cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1233 qb4 clk a_108_n1569# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1234 a_110_n119# a_55_n115# gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1235 q1 a_243_n281# p1 Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1236 g1_bar q6 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1237 q6 qb6 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1238 a_848_n913# g2 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 c4 a_849_n1172# vdd vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1240 a_875_n1667# g0 gnd Gnd cmosn w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1241 q4 a_240_n1589# p4 Gnd cmosn w=10 l=2
+  ad=100 pd=60 as=0 ps=0
M1242 a_871_n225# g0 gnd Gnd cmosn w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1243 a_838_n1779# p4 a_871_n1747# Gnd cmosn w=60 l=2
+  ad=300 pd=130 as=0 ps=0
M1244 a_47_n256# clk gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1245 c2 a_832_n299# vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1246 a_17_n585# a2 gnd Gnd cmosn w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1247 g3_bar q8 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1248 a_53_n1216# a_15_n1216# a_45_n1216# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1249 a_15_n1706# b4 gnd Gnd cmosn w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1250 a_19_23# clk a_19_46# vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1251 qb2 clk a_110_n589# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1252 a_55_n727# a_17_n727# a_47_n704# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1253 g3_bar a_225_n1179# a_279_n1185# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1254 a_243_n281# q6 vdd vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1255 c3 a_840_n663# vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 a_873_n647# p1 a_873_n655# Gnd cmosn w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1257 vdd p1 a_842_n1077# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1258 a_1098_n1540# a_841_n1482# a_1098_n1548# Gnd cmosn w=60 l=2
+  ad=0 pd=0 as=0 ps=0
M1259 q3 qb3 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1260 a_15_n2012# c0 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1261 a_55_n1075# a_17_n1075# a_47_n1075# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1262 a_875_n1061# p2 a_875_n1069# Gnd cmosn w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1263 a_15_n1193# b3 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1264 a_108_n1710# a_53_n1706# gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1265 a_112_19# a_57_23# gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1266 a_874_36# qc0 gnd Gnd cmosn w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1267 vdd p3 a_848_n1667# vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1268 a_840_n573# p2 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1269 a_873_n565# p1 a_873_n573# Gnd cmosn w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M1270 a_17_n375# b1 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1271 g3 g3_bar vdd vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1272 vdd p0 a_849_n1172# vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1273 a_847_n1408# g3 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1274 vdd q4 g4_bar vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1275 q9 qb9 vdd vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1276 g0_bar q0 a_281_n84# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1277 a_875_n987# g1 gnd Gnd cmosn w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M1278 c2 a_838_n225# a_1057_n246# Gnd cmosn w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M1279 a_1066_n577# a_840_n573# a_1066_n585# Gnd cmosn w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1280 qbc0 a_53_n2035# vdd vdd cmosp w=20 l=2
+  ad=260 pd=66 as=0 ps=0
M1281 a_838_n1779# qc0 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1282 a_57_23# a_19_23# a_49_23# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1283 a_832_n299# p1 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1284 a_865_n291# p0 a_865_n299# Gnd cmosn w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M1285 a_47_n398# clk gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1286 a_848_n913# p3 a_881_n913# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1287 c4 g3_bar vdd vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1288 a_53_n1706# a_15_n1706# a_45_n1706# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1289 q4 qb4 gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1290 q2 qb2 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1291 a_17_n1052# a3 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1292 a_875_n1651# p2 a_875_n1659# Gnd cmosn w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1293 a_876_n1172# qc0 gnd Gnd cmosn w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1294 a_871_n1763# p1 a_871_n1771# Gnd cmosn w=60 l=2
+  ad=0 pd=0 as=0 ps=0
M1295 a_15_n1565# clk a_15_n1542# vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1296 a_53_n2035# a_15_n2035# a_45_n2012# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1297 vdd q0 g0_bar vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1298 a_53_n1216# a_15_n1216# a_45_n1193# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1299 cout a_838_n1779# vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1300 a_841_n1572# g1 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1301 a_17_n727# b2 gnd Gnd cmosn w=10 l=2
+  ad=130 pd=46 as=0 ps=0
M1302 a_15_n1683# b4 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1303 a_240_n1589# q9 gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1304 a_847_n1408# p4 a_880_n1408# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1305 vdd p2 a_838_n1779# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1306 a_1098_n1564# a_848_n1667# a_1098_n1572# Gnd cmosn w=60 l=2
+  ad=0 pd=0 as=0 ps=0
M1307 a_874_n1564# p2 a_874_n1572# Gnd cmosn w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1308 p0 q0 a_243_2# Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1309 p1 q1 a_243_n281# Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1310 p4 q4 q9 vdd cmosp w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1311 a_17_n92# b0 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1312 a_848_n1667# g0 vdd vdd cmosp w=14 l=2
+  ad=0 pd=0 as=0 ps=0
M1313 g0 g0_bar gnd Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1314 a_874_n1482# g2 gnd Gnd cmosn w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M1315 qb5 a_55_n115# vdd vdd cmosp w=20 l=2
+  ad=260 pd=66 as=0 ps=0
M1316 a_47_n233# clk vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1317 a_17_n562# a2 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1318 qb1 a_55_n256# vdd vdd cmosp w=20 l=2
+  ad=260 pd=66 as=0 ps=0
M1319 a_876_n1148# p2 a_876_n1156# Gnd cmosn w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1320 a_842_n987# p3 a_875_n979# Gnd cmosn w=30 l=2
+  ad=150 pd=70 as=0 ps=0
M1321 vdd p1 a_838_n225# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1322 q2 a_243_n610# p2 Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1323 g2_bar q7 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1324 qbc0 clk a_108_n2039# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1325 a_57_23# a_19_23# a_49_46# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1326 vdd g4_bar cout vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1327 vdd p4 a_841_n1572# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1328 a_243_n281# q6 gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1329 a_846_n499# g1 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1330 a_55_n1075# a_17_n1075# a_47_n1052# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1331 a_45_n1565# clk gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1332 vdd p0 a_841_36# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1333 q1 q6 p1 vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1334 a_55_n115# rst vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1335 a_47_n585# clk gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1336 a_53_n1565# a_83_n1543# vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1337 a_55_n398# rst vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1338 a_841_n1482# p4 vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1339 q4 q9 p4 vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1340 c4 a_848_n913# a_1091_n1032# Gnd cmosn w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1341 a_243_n610# q7 vdd vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1342 a_53_n1706# a_15_n1706# a_45_n1683# vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_241_n1099# vdd 0.25fF
C1 a_840_n663# a_873_n655# 0.05fF
C2 p2 a_848_n1667# 0.08fF
C3 clk a_55_n585# 0.03fF
C4 a_53_n1216# a_15_n1216# 0.01fF
C5 a_842_n1077# a_849_n1172# 0.56fF
C6 a_1066_n593# gnd 0.41fF
C7 a1 clk 0.10fF
C8 g2_bar vdd 0.97fF
C9 a_875_n1643# a_848_n1667# 0.57fF
C10 a_847_n1408# a_880_n1408# 0.26fF
C11 vdd qbc0 0.41fF
C12 p4 g0_bar 0.14fF
C13 vdd g4_bar 0.98fF
C14 p2 a_840_n573# 0.08fF
C15 a0 clk 0.10fF
C16 a_838_n1779# a_871_n1771# 0.05fF
C17 a_17_n398# clk 0.27fF
C18 a_55_n398# rst 0.06fF
C19 a_17_n727# gnd 0.10fF
C20 g3_bar g4 0.16fF
C21 qb0 gnd 0.05fF
C22 a_846_n499# c3 0.08fF
C23 a_17_n398# a_17_n375# 0.21fF
C24 a_840_n663# p1 0.08fF
C25 gnd qc0 0.41fF
C26 a_874_n1556# a_874_n1564# 0.41fF
C27 p1 p4 0.47fF
C28 a_841_36# g0_bar 0.26fF
C29 a_47_n727# gnd 0.10fF
C30 g2_bar g3_bar 0.15fF
C31 g1_bar p4 0.16fF
C32 qb7 vdd 0.41fF
C33 a_1066_n585# a_1066_n577# 0.41fF
C34 a_875_n987# gnd 0.31fF
C35 q0 gnd 0.21fF
C36 p3 qc0 0.33fF
C37 p2 g4 0.52fF
C38 a_45_n1706# gnd 0.10fF
C39 g3_bar g4_bar 0.16fF
C40 qb3 gnd 0.05fF
C41 g3 p0 0.33fF
C42 qb8 gnd 0.05fF
C43 vdd g0_bar 0.97fF
C44 a_874_n1572# gnd 0.41fF
C45 a_110_n260# gnd 0.10fF
C46 a_847_n1408# cout 0.08fF
C47 clk qbc0 0.01fF
C48 a_848_n913# vdd 0.67fF
C49 g2_bar p2 0.52fF
C50 a_17_n115# gnd 0.10fF
C51 a3 vdd 0.19fF
C52 qb4 gnd 0.05fF
C53 p1 vdd 2.31fF
C54 a_281_n84# gnd 0.21fF
C55 a_17_n115# a_55_n115# 0.01fF
C56 a_17_n1075# a_17_n1052# 0.21fF
C57 a_15_n1216# a_15_n1193# 0.21fF
C58 p2 g4_bar 0.61fF
C59 gnd a_17_n585# 0.10fF
C60 a_1057_n254# gnd 0.31fF
C61 g1_bar vdd 0.99fF
C62 gnd a_110_n589# 0.10fF
C63 a_838_n225# a_871_n225# 0.26fF
C64 c4 vdd 0.88fF
C65 vdd a_15_n1565# 0.77fF
C66 qb5 vdd 0.41fF
C67 g3_bar g0_bar 0.14fF
C68 q8 qb8 0.05fF
C69 c4 a_1091_n1056# 0.05fF
C70 qb7 clk 0.01fF
C71 a_19_23# gnd 0.10fF
C72 q5 a_243_2# 0.05fF
C73 q1 vdd 1.05fF
C74 c0 a_15_n2012# 0.01fF
C75 a_53_n2035# a_45_n2012# 0.21fF
C76 vdd qb2 0.41fF
C77 p1 a_832_n299# 0.08fF
C78 g0 a_848_n1667# 0.08fF
C79 p4 a_841_n1572# 0.08fF
C80 g1 qc0 0.33fF
C81 p1 g3_bar 0.47fF
C82 g1_bar a_832_n299# 0.31fF
C83 g2 g4 0.19fF
C84 c2 a_1057_n254# 0.05fF
C85 a_841_n1572# a_874_n1556# 0.47fF
C86 p2 g0_bar 0.14fF
C87 a_849_n1172# a_876_n1148# 0.57fF
C88 a_55_n398# vdd 0.80fF
C89 g1_bar g3_bar 0.16fF
C90 rst a_57_23# 0.06fF
C91 a3 clk 0.10fF
C92 a_53_n1216# gnd 0.05fF
C93 a_1098_n1564# cout 0.05fF
C94 c4 g3_bar 0.08fF
C95 q3 a_225_n1179# 0.03fF
C96 g2_bar g2 22.62fF
C97 a_842_n1077# a_875_n1061# 0.47fF
C98 vdd a_45_n1683# 0.21fF
C99 a_53_n2035# gnd 0.05fF
C100 p1 p2 5.61fF
C101 clk a_15_n1565# 0.27fF
C102 rst a_53_n1565# 0.05fF
C103 a_108_n2039# gnd 0.10fF
C104 qb5 clk 0.01fF
C105 g1_bar p2 22.33fF
C106 g2 g4_bar 0.19fF
C107 q4 qb4 0.05fF
C108 a_840_n573# c3 0.08fF
C109 a_840_n663# p0 0.08fF
C110 vdd a_841_n1572# 1.25fF
C111 a_838_n1779# a_871_n1763# 0.05fF
C112 clk qb2 0.01fF
C113 p3 a_842_n1077# 0.08fF
C114 c3 a_1066_n577# 0.47fF
C115 p4 p0 0.33fF
C116 vdd a_15_n2012# 0.21fF
C117 a_841_n1482# g4_bar 0.60fF
C118 g0 g4 0.28fF
C119 m4_437_29# qc0 0.05fF
C120 b2 a_17_n704# 0.01fF
C121 a_55_n398# clk 0.03fF
C122 a_873_n663# gnd 0.41fF
C123 a_19_23# a_19_46# 0.21fF
C124 a_281_n696# gnd 0.21fF
C125 gnd a_243_2# 0.10fF
C126 p0 a_841_36# 0.08fF
C127 g2_bar g0 0.28fF
C128 g3_bar a_279_n1185# 0.26fF
C129 a_875_n1667# gnd 0.52fF
C130 g2 g0_bar 0.14fF
C131 a_841_36# a_874_36# 0.26fF
C132 g3 p4 0.95fF
C133 g0 g4_bar 0.28fF
C134 a_17_n704# vdd 0.21fF
C135 a_871_n1763# a_871_n1771# 0.62fF
C136 g2_bar c3 0.08fF
C137 vdd p0 1.49fF
C138 b4 a_15_n1683# 0.01fF
C139 a_57_23# a_49_46# 0.21fF
C140 q0 qb0 0.05fF
C141 a_53_n1706# a_45_n1683# 0.21fF
C142 g2 p1 0.47fF
C143 p4 q9 0.29fF
C144 a_871_n225# gnd 0.21fF
C145 g2 g1_bar 0.16fF
C146 a_848_n913# a_881_n913# 0.26fF
C147 p3 a_842_n987# 0.08fF
C148 p2 a_841_n1572# 0.08fF
C149 a_848_n1667# gnd 0.18fF
C150 a_1091_n1040# a_1091_n1048# 0.52fF
C151 p1 a_849_n1172# 0.08fF
C152 q3 vdd 0.84fF
C153 vdd a_57_23# 0.80fF
C154 qb1 vdd 0.41fF
C155 g3 vdd 0.62fF
C156 gnd a_55_n585# 0.05fF
C157 a_832_n299# p0 0.08fF
C158 p3 a_848_n1667# 0.08fF
C159 a_243_n281# vdd 0.25fF
C160 g0 g0_bar 22.67fF
C161 qb7 q7 0.05fF
C162 p1 a_838_n225# 0.08fF
C163 g3_bar p0 0.33fF
C164 vdd a_53_n1565# 0.80fF
C165 a_17_n92# vdd 0.21fF
C166 a_838_n225# g1_bar 0.31fF
C167 vdd q9 1.38fF
C168 a_53_n2035# a_15_n2035# 0.01fF
C169 p1 g0 3.26fF
C170 vdd a_17_n562# 0.21fF
C171 a_17_n398# gnd 0.10fF
C172 vdd a_243_n610# 0.25fF
C173 p2 p0 0.33fF
C174 a_110_n402# gnd 0.10fF
C175 g1_bar g0 0.28fF
C176 c4 a_1091_n1032# 0.57fF
C177 a_874_n1474# a_874_n1482# 0.31fF
C178 a_838_n1779# a_848_n1667# 0.28fF
C179 cout a_848_n1667# 0.08fF
C180 g3_bar g3 22.36fF
C181 g4 gnd 0.10fF
C182 a_53_n1565# a_45_n1542# 0.21fF
C183 a4 a_15_n1542# 0.01fF
C184 rst vdd 5.54fF
C185 clk a_57_23# 0.03fF
C186 a_241_n1099# gnd 0.10fF
C187 qb1 clk 0.01fF
C188 qb6 vdd 0.41fF
C189 a_225_n1179# vdd 0.20fF
C190 a_55_n585# a_47_n562# 0.21fF
C191 a2 a_17_n562# 0.01fF
C192 p3 g4 0.47fF
C193 g2_bar gnd 0.24fF
C194 vdd a_15_n1706# 0.77fF
C195 a_838_n1779# a_871_n1755# 0.05fF
C196 a_876_n1148# a_876_n1156# 0.52fF
C197 p3 a_241_n1099# 0.20fF
C198 clk a_53_n1565# 0.03fF
C199 p2 g3 0.52fF
C200 a_45_n1216# gnd 0.10fF
C201 qb5 q5 0.05fF
C202 qbc0 gnd 0.05fF
C203 b3 vdd 0.19fF
C204 q9 a_240_n1589# 0.05fF
C205 g4_bar gnd 22.39fF
C206 a_840_n573# a_873_n565# 0.36fF
C207 g2_bar p3 22.31fF
C208 a_1098_n1548# a_1098_n1556# 0.62fF
C209 vdd c0 0.19fF
C210 a_873_n647# a_873_n655# 0.41fF
C211 q8 a_241_n1099# 0.05fF
C212 p3 g4_bar 0.47fF
C213 g3_bar a_225_n1179# 0.08fF
C214 p2 a_243_n610# 0.20fF
C215 a0 a_19_46# 0.01fF
C216 a_840_n663# vdd 1.21fF
C217 clk rst 0.55fF
C218 qb6 clk 0.01fF
C219 qb7 gnd 0.05fF
C220 g2 p0 0.33fF
C221 gnd a_49_23# 0.10fF
C222 p4 vdd 1.40fF
C223 a_55_n398# a_47_n398# 0.10fF
C224 clk a_15_n1706# 0.27fF
C225 rst a_53_n1706# 0.06fF
C226 gnd g0_bar 0.20fF
C227 a_849_n1172# p0 0.08fF
C228 b2 vdd 0.19fF
C229 b3 clk 0.10fF
C230 g1 g4 0.24fF
C231 vdd a_49_46# 0.21fF
C232 cout g4_bar 0.08fF
C233 a_53_n1706# a_15_n1706# 0.01fF
C234 p3 g0_bar 0.14fF
C235 vdd a_841_36# 0.71fF
C236 q0 a_243_2# 0.01fF
C237 g2 g3 0.19fF
C238 p1 gnd 0.37fF
C239 clk c0 0.10fF
C240 p3 a_848_n913# 0.08fF
C241 g1_bar gnd 0.23fF
C242 g2_bar g1 0.24fF
C243 a_842_n987# a_875_n987# 0.05fF
C244 g3_bar p4 22.33fF
C245 q4 g4_bar 0.08fF
C246 g2_bar q2 0.08fF
C247 p1 p3 0.48fF
C248 a_15_n1565# gnd 0.10fF
C249 qb5 gnd 0.05fF
C250 g0 p0 22.55fF
C251 a_875_n1643# a_875_n1651# 0.52fF
C252 a_47_n1052# vdd 0.21fF
C253 a_45_n1193# vdd 0.21fF
C254 g1 g4_bar 0.24fF
C255 a_45_n1565# gnd 0.10fF
C256 p4 a_240_n1589# 0.20fF
C257 g1_bar p3 0.16fF
C258 q1 gnd 0.20fF
C259 a_17_n92# b0 0.01fF
C260 gnd qb2 0.05fF
C261 a_1098_n1540# a_1098_n1548# 0.62fF
C262 q6 p1 0.29fF
C263 a_840_n663# p2 0.08fF
C264 a_875_n1077# gnd 0.41fF
C265 gnd a_873_n573# 0.31fF
C266 p2 p4 0.52fF
C267 b2 clk 0.10fF
C268 a_55_n727# rst 0.06fF
C269 a_841_n1482# a_874_n1482# 0.05fF
C270 q5 p0 0.29fF
C271 vdd a_45_n1542# 0.21fF
C272 c2 g1_bar 0.08fF
C273 vdd a2 0.19fF
C274 a_55_n398# gnd 0.05fF
C275 a_832_n299# vdd 0.96fF
C276 g0 g3 0.28fF
C277 a_17_n256# vdd 0.77fF
C278 a_110_n1079# gnd 0.10fF
C279 p1 a_838_n1779# 0.08fF
C280 g3_bar vdd 1.02fF
C281 q6 q1 0.88fF
C282 a_281_n367# gnd 0.21fF
C283 a_53_n1565# a_83_n1543# 0.01fF
C284 g1 g0_bar 0.14fF
C285 vdd a_240_n1589# 0.25fF
C286 a_838_n1779# a_871_n1747# 0.67fF
C287 clk vdd 11.44fF
C288 g4 qc0 0.33fF
C289 qb5 a_110_n119# 0.10fF
C290 a_17_n375# vdd 0.21fF
C291 a_279_n1185# gnd 0.21fF
C292 a_841_n1572# gnd 0.18fF
C293 p2 vdd 2.58fF
C294 vdd a_53_n1706# 0.80fF
C295 a_55_n585# a_17_n585# 0.01fF
C296 p1 g1 22.77fF
C297 g2_bar qc0 0.33fF
C298 a1 a_17_n233# 0.01fF
C299 qb9 a_108_n1710# 0.10fF
C300 g1_bar g1 22.61fF
C301 q7 a_243_n610# 0.05fF
C302 rst a_83_n1543# 0.05fF
C303 p3 a_841_n1572# 0.08fF
C304 qbc0 qc0 0.05fF
C305 clk a2 0.10fF
C306 a_278_n1675# gnd 0.21fF
C307 g4_bar qc0 0.33fF
C308 a_873_n565# a_873_n573# 0.31fF
C309 a_55_n256# rst 0.06fF
C310 a_17_n256# clk 0.27fF
C311 g2 p4 0.19fF
C312 a_871_n1755# a_871_n1763# 0.62fF
C313 qb9 q9 0.05fF
C314 p2 g3_bar 0.52fF
C315 q2 qb2 0.05fF
C316 a_846_n499# a_840_n573# 0.37fF
C317 p4 a_841_n1482# 0.08fF
C318 p0 gnd 0.23fF
C319 cout a_841_n1572# 0.08fF
C320 clk a_53_n1706# 0.03fF
C321 gnd a_874_36# 0.21fF
C322 qc0 g0_bar 0.33fF
C323 a_55_n727# vdd 0.80fF
C324 p3 p0 0.33fF
C325 a_110_n731# gnd 0.10fF
C326 g1_bar m4_437_29# 0.00fF
C327 c4 a_1091_n1048# 0.05fF
C328 g2 vdd 0.89fF
C329 q3 gnd 0.28fF
C330 a_57_23# gnd 0.05fF
C331 a_108_n1710# gnd 0.10fF
C332 qb1 gnd 0.05fF
C333 g3 gnd 0.15fF
C334 g0 p4 0.28fF
C335 q0 g0_bar 0.08fF
C336 vdd b0 0.19fF
C337 g1 a_841_n1572# 0.08fF
C338 a_849_n1172# vdd 1.12fF
C339 a_243_n281# gnd 0.10fF
C340 p1 qc0 0.32fF
C341 p3 q3 0.51fF
C342 a_841_n1482# vdd 0.96fF
C343 a_875_n1061# a_875_n1069# 0.41fF
C344 g1_bar qc0 0.33fF
C345 a_53_n1565# gnd 0.05fF
C346 a_875_n1667# a_848_n1667# 0.05fF
C347 p3 g3 22.75fF
C348 a_15_n1216# vdd 0.77fF
C349 a_17_n1075# vdd 0.77fF
C350 a_838_n1779# p0 0.08fF
C351 q9 gnd 0.25fF
C352 a_47_n115# gnd 0.10fF
C353 a_838_n225# vdd 0.63fF
C354 a_841_n1482# a_874_n1474# 0.36fF
C355 a_874_n1482# gnd 0.31fF
C356 cout a_1098_n1556# 0.05fF
C357 a_874_n1572# a_874_n1564# 0.41fF
C358 a_281_n84# g0_bar 0.26fF
C359 a_47_n115# a_55_n115# 0.10fF
C360 g2 g3_bar 0.19fF
C361 q6 a_243_n281# 0.05fF
C362 a_53_n1216# a_45_n1216# 0.10fF
C363 gnd a_243_n610# 0.10fF
C364 q3 q8 0.58fF
C365 a_55_n727# clk 0.03fF
C366 vdd a_83_n1543# 0.21fF
C367 g0 vdd 1.49fF
C368 rst gnd 0.54fF
C369 a_55_n256# vdd 0.80fF
C370 a_15_n2035# a_15_n2012# 0.21fF
C371 a_849_n1172# a_876_n1172# 0.05fF
C372 g1 p0 0.33fF
C373 qb6 gnd 0.05fF
C374 vdd q7 1.46fF
C375 clk b0 0.10fF
C376 rst a_55_n115# 0.06fF
C377 qbc0 a_108_n2039# 0.10fF
C378 g2 p2 22.81fF
C379 vdd c3 1.01fF
C380 a_47_n256# a_55_n256# 0.10fF
C381 a_879_n499# gnd 0.21fF
C382 a_15_n1706# gnd 0.10fF
C383 q5 vdd 1.39fF
C384 p2 a_849_n1172# 0.08fF
C385 b1 vdd 0.19fF
C386 a_55_n1075# rst 0.06fF
C387 a_17_n1075# clk 0.27fF
C388 a_15_n1216# clk 0.27fF
C389 c4 a_1091_n1040# 0.05fF
C390 qb3 a_110_n1079# 0.10fF
C391 q6 qb6 0.05fF
C392 g0 g3_bar 0.28fF
C393 g2_bar a_281_n696# 0.26fF
C394 g1 g3 0.24fF
C395 a_55_n256# a_17_n256# 0.01fF
C396 vdd qb9 0.41fF
C397 a_876_n1164# a_876_n1172# 0.52fF
C398 a_840_n663# a_873_n647# 0.47fF
C399 qb2 a_110_n589# 0.10fF
C400 q8 a_225_n1179# 0.26fF
C401 q4 q9 0.78fF
C402 a_55_n256# clk 0.03fF
C403 g0 p2 0.28fF
C404 p4 gnd 0.23fF
C405 vdd a_45_n2012# 0.21fF
C406 a_874_n1572# a_841_n1572# 0.05fF
C407 cout a_1098_n1540# 0.67fF
C408 a_873_n655# a_873_n663# 0.41fF
C409 p1 a_842_n1077# 0.08fF
C410 p2 q7 0.29fF
C411 a_17_n727# a_17_n704# 0.21fF
C412 b1 clk 0.10fF
C413 q2 a_243_n610# 0.01fF
C414 a_875_n1659# a_875_n1667# 0.52fF
C415 p3 p4 3.66fF
C416 a_55_n398# a_47_n375# 0.21fF
C417 b1 a_17_n375# 0.01fF
C418 c4 a_842_n1077# 0.08fF
C419 p0 qc0 26.58fF
C420 gnd a_841_36# 0.06fF
C421 a_832_n299# a_865_n299# 0.05fF
C422 clk qb9 0.01fF
C423 g2_bar a_840_n573# 0.60fF
C424 a_47_n704# vdd 0.21fF
C425 a_1066_n585# c3 0.05fF
C426 vdd gnd 7.07fF
C427 a_15_n1706# a_15_n1683# 0.21fF
C428 q0 p0 0.51fF
C429 a_842_n1077# a_875_n1077# 0.05fF
C430 vdd a_55_n115# 0.80fF
C431 a_1091_n1056# gnd 0.52fF
C432 a_875_n1659# a_848_n1667# 0.05fF
C433 p4 a_838_n1779# 0.08fF
C434 a_47_n256# gnd 0.10fF
C435 g3 qc0 0.33fF
C436 a_848_n913# a_842_n987# 0.40fF
C437 p3 vdd 2.23fF
C438 a_55_n1075# vdd 0.80fF
C439 g2_bar g4 0.15fF
C440 g2 g0 0.28fF
C441 q6 vdd 1.39fF
C442 a_970_n61# gnd 0.21fF
C443 a_55_n1075# a_47_n1052# 0.21fF
C444 q3 qb3 0.05fF
C445 a3 a_17_n1052# 0.01fF
C446 a_1098_n1564# a_1098_n1556# 0.62fF
C447 p4 q4 0.51fF
C448 c2 vdd 0.76fF
C449 a_17_n256# gnd 0.10fF
C450 gnd a_47_n585# 0.10fF
C451 a_849_n1172# a_876_n1164# 0.05fF
C452 g4 g4_bar 22.29fF
C453 g3_bar gnd 0.25fF
C454 qb1 a_110_n260# 0.10fF
C455 a_842_n987# c4 0.08fF
C456 g1 p4 0.25fF
C457 q8 vdd 1.40fF
C458 vdd a4 0.19fF
C459 a_876_n1172# gnd 0.52fF
C460 a_47_n92# vdd 0.21fF
C461 p1 a_848_n1667# 0.08fF
C462 a_240_n1589# gnd 0.10fF
C463 vdd a_838_n1779# 1.72fF
C464 vdd cout 1.52fF
C465 clk gnd 11.29fF
C466 p3 g3_bar 0.47fF
C467 g2_bar g4_bar 0.15fF
C468 vdd a_47_n562# 0.21fF
C469 clk a_55_n115# 0.03fF
C470 p2 gnd 0.42fF
C471 a_53_n1706# gnd 0.05fF
C472 p1 a_840_n573# 0.08fF
C473 a_17_n115# a_17_n92# 0.21fF
C474 a_15_n1565# a_15_n1542# 0.21fF
C475 vdd q4 1.06fF
C476 a_55_n1075# clk 0.03fF
C477 a_19_23# a_57_23# 0.01fF
C478 a_19_46# vdd 0.21fF
C479 g4 g0_bar 0.14fF
C480 p2 p3 5.47fF
C481 g1 vdd 1.17fF
C482 a_871_n1747# a_871_n1755# 0.62fF
C483 q2 vdd 1.05fF
C484 a_17_n585# a_17_n562# 0.21fF
C485 vdd a_15_n1683# 0.21fF
C486 clk a4 0.10fF
C487 g2_bar g0_bar 0.14fF
C488 p4 a_847_n1408# 0.08fF
C489 a_45_n2035# gnd 0.10fF
C490 a_108_n1220# gnd 0.10fF
C491 p1 g4 0.47fF
C492 a_840_n573# a_873_n573# 0.05fF
C493 a_832_n299# a_865_n291# 0.36fF
C494 g1_bar g4 0.16fF
C495 g4_bar g0_bar 0.14fF
C496 p2 a_838_n1779# 0.08fF
C497 vdd a_15_n2035# 0.77fF
C498 g2_bar p1 0.47fF
C499 p4 qc0 0.33fF
C500 g1 g3_bar 0.24fF
C501 a_841_n1572# a_848_n1667# 0.45fF
C502 q4 a_240_n1589# 0.01fF
C503 a_55_n727# a_47_n704# 0.21fF
C504 g2_bar g1_bar 0.16fF
C505 a_55_n727# gnd 0.05fF
C506 p1 g4_bar 0.47fF
C507 a_55_n398# a_17_n398# 0.01fF
C508 g2 gnd 0.20fF
C509 gnd a_112_19# 0.10fF
C510 p0 a_243_2# 0.19fF
C511 a_847_n1408# vdd 0.71fF
C512 g1_bar g4_bar 0.16fF
C513 a_842_n1077# a_875_n1069# 0.05fF
C514 a_1091_n1048# a_1091_n1056# 0.52fF
C515 g1 p2 2.75fF
C516 a_849_n1172# gnd 0.06fF
C517 g2 p3 1.86fF
C518 a_17_n727# vdd 0.77fF
C519 a_881_n913# gnd 0.21fF
C520 a_846_n499# a_879_n499# 0.26fF
C521 p2 q2 0.51fF
C522 vdd qb0 0.41fF
C523 a_53_n1216# rst 0.06fF
C524 cout a_1098_n1548# 0.05fF
C525 a_15_n1216# gnd 0.10fF
C526 a_17_n1075# gnd 0.10fF
C527 vdd qc0 1.70fF
C528 p3 a_849_n1172# 0.08fF
C529 p3 a_841_n1482# 0.08fF
C530 rst a_53_n2035# 0.01fF
C531 clk a_15_n2035# 0.27fF
C532 p1 g0_bar 22.29fF
C533 a_849_n1172# a_876_n1156# 0.05fF
C534 a_875_n979# a_875_n987# 0.31fF
C535 vdd q0 1.06fF
C536 g1_bar g0_bar 0.14fF
C537 g0 gnd 0.29fF
C538 a_47_n233# vdd 0.21fF
C539 a_55_n1075# a_17_n1075# 0.01fF
C540 qb3 vdd 0.41fF
C541 qb8 vdd 0.41fF
C542 a_108_n1569# gnd 0.10fF
C543 a_55_n256# gnd 0.05fF
C544 gnd q7 0.27fF
C545 a_848_n913# c4 0.08fF
C546 g0 p3 0.28fF
C547 a_17_n115# vdd 0.77fF
C548 a_838_n225# c2 0.08fF
C549 p1 g1_bar 0.47fF
C550 g3_bar qc0 0.33fF
C551 a_1098_n1572# gnd 0.62fF
C552 a_841_n1482# cout 0.08fF
C553 a_17_n727# clk 0.27fF
C554 clk qb0 0.01fF
C555 q5 gnd 0.27fF
C556 vdd qb4 0.41fF
C557 c2 a_1057_n246# 0.36fF
C558 a_841_n1572# g4_bar 0.61fF
C559 vdd a_17_n585# 0.77fF
C560 a_876_n1156# a_876_n1164# 0.52fF
C561 a_17_n233# vdd 0.21fF
C562 g2 g1 0.24fF
C563 p1 q1 0.51fF
C564 a_1066_n585# a_1066_n593# 0.41fF
C565 a_47_n398# gnd 0.10fF
C566 p2 qc0 0.33fF
C567 g1_bar q1 0.08fF
C568 qb9 gnd 0.05fF
C569 g4 p0 0.33fF
C570 a_19_23# vdd 0.77fF
C571 a_278_n1675# g4_bar 0.26fF
C572 a_47_n375# vdd 0.21fF
C573 qb3 clk 0.01fF
C574 qb8 clk 0.01fF
C575 a_865_n299# gnd 0.31fF
C576 a_846_n499# vdd 0.71fF
C577 g2_bar p0 0.33fF
C578 vdd b4 0.19fF
C579 a_53_n1706# a_45_n1706# 0.10fF
C580 a_871_n1779# gnd 0.62fF
C581 a_17_n256# a_17_n233# 0.21fF
C582 a_17_n115# clk 0.27fF
C583 g1_bar a_281_n367# 0.26fF
C584 a_53_n1216# vdd 0.80fF
C585 a_1098_n1572# cout 0.05fF
C586 q3 a_241_n1099# 0.01fF
C587 a_840_n663# a_873_n663# 0.05fF
C588 clk qb4 0.01fF
C589 g3 g4 0.14fF
C590 g4_bar p0 0.33fF
C591 b3 a_15_n1193# 0.01fF
C592 a_841_n1572# a_874_n1564# 0.05fF
C593 a_53_n1216# a_45_n1193# 0.21fF
C594 rst a_55_n585# 0.06fF
C595 clk a_17_n585# 0.27fF
C596 g0 g1 0.28fF
C597 vdd a_53_n2035# 0.80fF
C598 a_842_n1077# vdd 1.25fF
C599 g2_bar g3 0.15fF
C600 a_55_n727# a_17_n727# 0.01fF
C601 q2 q7 0.83fF
C602 clk a_19_23# 0.27fF
C603 qb8 a_108_n1220# 0.10fF
C604 a_875_n1651# a_848_n1667# 0.05fF
C605 g3 g4_bar 0.14fF
C606 a_847_n1408# a_841_n1482# 0.36fF
C607 qb0 a_112_19# 0.10fF
C608 a_880_n1408# gnd 0.21fF
C609 clk b4 0.10fF
C610 g2 qc0 0.33fF
C611 a_55_n727# a_47_n727# 0.10fF
C612 p0 g0_bar 0.33fF
C613 gnd a_55_n115# 0.05fF
C614 a_838_n1779# a_871_n1779# 0.05fF
C615 qb6 a_110_n402# 0.10fF
C616 qb7 a_110_n731# 0.10fF
C617 p2 a_846_n499# 0.08fF
C618 p3 gnd 0.37fF
C619 a_53_n1216# clk 0.03fF
C620 g3_bar a_842_n1077# 0.93fF
C621 p4 a_848_n1667# 0.08fF
C622 a_55_n1075# gnd 0.05fF
C623 a_57_23# a_49_23# 0.10fF
C624 vdd a_243_2# 0.25fF
C625 a_865_n291# a_865_n299# 0.31fF
C626 q6 gnd 0.27fF
C627 p1 p0 3.93fF
C628 clk a_53_n2035# 0.03fF
C629 g1_bar p0 0.33fF
C630 g3 g0_bar 0.14fF
C631 a_1066_n593# c3 0.05fF
C632 a_842_n987# a_875_n979# 0.36fF
C633 q8 gnd 0.27fF
C634 a_842_n987# vdd 1.00fF
C635 p2 a_842_n1077# 0.08fF
C636 a_17_n1052# vdd 0.21fF
C637 a_15_n1193# vdd 0.21fF
C638 a_838_n1779# gnd 0.06fF
C639 g0 qc0 0.32fF
C640 a_871_n1771# a_871_n1779# 0.62fF
C641 c1 a_841_36# 0.08fF
C642 a_47_n92# a_55_n115# 0.21fF
C643 a_110_n119# gnd 0.10fF
C644 p3 q8 0.29fF
C645 p1 g3 0.47fF
C646 vdd a_848_n1667# 1.12fF
C647 p1 a_243_n281# 0.19fF
C648 g1_bar g3 0.16fF
C649 p3 a_838_n1779# 0.08fF
C650 vdd a_15_n1542# 0.21fF
C651 c1 vdd 0.51fF
C652 p4 g4 22.56fF
C653 vdd a_55_n585# 0.80fF
C654 q4 gnd 0.30fF
C655 a1 vdd 0.19fF
C656 a_53_n2035# a_45_n2035# 0.10fF
C657 a_47_n1075# gnd 0.10fF
C658 vdd a_840_n573# 0.96fF
C659 a_842_n987# g3_bar 0.71fF
C660 g2_bar a_840_n663# 0.37fF
C661 g1 gnd 0.24fF
C662 qb1 q1 0.05fF
C663 a_47_n233# a_55_n256# 0.21fF
C664 a_243_n281# q1 0.01fF
C665 a_53_n1565# a_15_n1565# 0.01fF
C666 q2 gnd 0.30fF
C667 g2_bar p4 0.15fF
C668 q5 q0 0.78fF
C669 a_1057_n246# a_1057_n254# 0.31fF
C670 a0 vdd 0.19fF
C671 a_53_n1565# a_45_n1565# 0.10fF
C672 a_17_n398# vdd 0.77fF
C673 g1 p3 0.24fF
C674 c1 a_970_n61# 0.26fF
C675 a_875_n1651# a_875_n1659# 0.52fF
C676 a_55_n1075# a_47_n1075# 0.10fF
C677 qb4 a_108_n1569# 0.10fF
C678 p4 g4_bar 0.34fF
C679 p2 a_842_n987# 0.08fF
C680 a_1091_n1032# a_1091_n1040# 0.52fF
C681 a_875_n1069# a_875_n1077# 0.41fF
C682 a_55_n585# a_47_n585# 0.10fF
C683 vdd g4 0.35fF
C684 a_15_n2035# gnd 0.10fF
C685 a_1098_n1564# a_1098_n1572# 0.62fF
C686 m4_437_29# Gnd 0.00fF 
C687 a_108_n2039# Gnd 0.01fF
C688 a_45_n2035# Gnd 0.01fF
C689 qbc0 Gnd 0.23fF
C690 a_15_n2035# Gnd 0.16fF
C691 c0 Gnd 0.08fF
C692 a_53_n2035# Gnd 0.23fF
C693 a_871_n1779# Gnd 0.01fF
C694 a_871_n1771# Gnd 0.01fF
C695 a_871_n1763# Gnd 0.01fF
C696 a_871_n1755# Gnd 0.01fF
C697 a_871_n1747# Gnd 0.01fF
C698 a_108_n1710# Gnd 0.01fF
C699 a_45_n1706# Gnd 0.01fF
C700 a_875_n1667# Gnd 0.01fF
C701 a_875_n1659# Gnd 0.01fF
C702 a_278_n1675# Gnd 0.01fF
C703 a_875_n1651# Gnd 0.01fF
C704 a_875_n1643# Gnd 0.01fF
C705 g4 Gnd 8.20fF
C706 qb9 Gnd 0.23fF
C707 a_15_n1706# Gnd 0.16fF
C708 b4 Gnd 0.08fF
C709 a_53_n1706# Gnd 0.23fF
C710 a_1098_n1572# Gnd 0.01fF
C711 a_838_n1779# Gnd 1.40fF
C712 a_874_n1572# Gnd 0.01fF
C713 a_1098_n1564# Gnd 0.01fF
C714 a_848_n1667# Gnd 1.39fF
C715 a_874_n1564# Gnd 0.01fF
C716 a_1098_n1556# Gnd 0.01fF
C717 a_874_n1556# Gnd 0.01fF
C718 a_1098_n1548# Gnd 0.01fF
C719 g4_bar Gnd 10.54fF
C720 a_841_n1572# Gnd 1.10fF
C721 a_1098_n1540# Gnd 0.01fF
C722 a_240_n1589# Gnd 0.41fF
C723 a_108_n1569# Gnd 0.01fF
C724 a_45_n1565# Gnd 0.01fF
C725 cout Gnd 0.18fF
C726 q9 Gnd 2.95fF
C727 qb4 Gnd 0.23fF
C728 a_83_n1543# Gnd 0.00fF
C729 a_15_n1565# Gnd 0.16fF
C730 a4 Gnd 0.08fF
C731 a_53_n1565# Gnd 0.23fF
C732 q4 Gnd 2.55fF
C733 a_874_n1482# Gnd 0.01fF
C734 a_874_n1474# Gnd 0.01fF
C735 a_841_n1482# Gnd 1.15fF
C736 a_880_n1408# Gnd 0.01fF
C737 a_847_n1408# Gnd 1.24fF
C738 p4 Gnd 12.29fF
C739 a_108_n1220# Gnd 0.01fF
C740 a_45_n1216# Gnd 0.01fF
C741 a_279_n1185# Gnd 0.01fF
C742 a_225_n1179# Gnd 0.17fF
C743 a_876_n1172# Gnd 0.01fF
C744 a_876_n1164# Gnd 0.01fF
C745 a_876_n1156# Gnd 0.01fF
C746 g3 Gnd 8.53fF
C747 qb8 Gnd 0.23fF
C748 a_15_n1216# Gnd 0.16fF
C749 b3 Gnd 0.08fF
C750 a_53_n1216# Gnd 0.23fF
C751 a_876_n1148# Gnd 0.01fF
C752 a_875_n1077# Gnd 0.01fF
C753 a_875_n1069# Gnd 0.01fF
C754 a_1091_n1056# Gnd 0.01fF
C755 a_849_n1172# Gnd 1.06fF
C756 a_875_n1061# Gnd 0.01fF
C757 a_1091_n1048# Gnd 0.01fF
C758 a_842_n1077# Gnd 0.84fF
C759 a_241_n1099# Gnd 0.41fF
C760 a_110_n1079# Gnd 0.01fF
C761 a_47_n1075# Gnd 0.01fF
C762 a_1091_n1040# Gnd 0.01fF
C763 g3_bar Gnd 10.50fF
C764 a_1091_n1032# Gnd 0.01fF
C765 c4 Gnd 0.15fF
C766 q8 Gnd 3.07fF
C767 qb3 Gnd 0.23fF
C768 a_17_n1075# Gnd 0.16fF
C769 a3 Gnd 0.08fF
C770 a_55_n1075# Gnd 0.23fF
C771 q3 Gnd 2.15fF
C772 a_875_n987# Gnd 0.01fF
C773 a_875_n979# Gnd 0.01fF
C774 a_842_n987# Gnd 1.08fF
C775 a_881_n913# Gnd 0.01fF
C776 a_848_n913# Gnd 1.17fF
C777 p3 Gnd 14.30fF
C778 a_110_n731# Gnd 0.01fF
C779 a_47_n727# Gnd 0.01fF
C780 a_281_n696# Gnd 0.01fF
C781 g2 Gnd 8.97fF
C782 qb7 Gnd 0.23fF
C783 a_17_n727# Gnd 0.16fF
C784 b2 Gnd 0.08fF
C785 a_873_n663# Gnd 0.01fF
C786 a_55_n727# Gnd 0.23fF
C787 a_873_n655# Gnd 0.01fF
C788 a_873_n647# Gnd 0.01fF
C789 a_1066_n593# Gnd 0.01fF
C790 a_840_n663# Gnd 0.84fF
C791 a_1066_n585# Gnd 0.01fF
C792 g2_bar Gnd 10.75fF
C793 a_1066_n577# Gnd 0.01fF
C794 c3 Gnd 0.13fF
C795 a_873_n573# Gnd 0.01fF
C796 a_873_n565# Gnd 0.01fF
C797 a_243_n610# Gnd 0.41fF
C798 a_110_n589# Gnd 0.01fF
C799 a_47_n585# Gnd 0.01fF
C800 a_840_n573# Gnd 0.85fF
C801 q7 Gnd 3.27fF
C802 qb2 Gnd 0.23fF
C803 a_17_n585# Gnd 0.16fF
C804 a2 Gnd 0.08fF
C805 a_55_n585# Gnd 0.23fF
C806 q2 Gnd 2.46fF
C807 a_879_n499# Gnd 0.01fF
C808 a_846_n499# Gnd 0.96fF
C809 p2 Gnd 14.36fF
C810 a_110_n402# Gnd 0.01fF
C811 a_47_n398# Gnd 0.01fF
C812 a_281_n367# Gnd 0.01fF
C813 g1 Gnd 9.47fF
C814 qb6 Gnd 0.23fF
C815 a_17_n398# Gnd 0.16fF
C816 b1 Gnd 0.08fF
C817 a_55_n398# Gnd 0.23fF
C818 a_865_n299# Gnd 0.01fF
C819 a_865_n291# Gnd 0.01fF
C820 a_1057_n254# Gnd 0.01fF
C821 a_832_n299# Gnd 0.76fF
C822 a_1057_n246# Gnd 0.01fF
C823 g1_bar Gnd 10.54fF
C824 c2 Gnd 0.11fF
C825 a_243_n281# Gnd 0.41fF
C826 a_110_n260# Gnd 0.01fF
C827 a_47_n256# Gnd 0.01fF
C828 a_871_n225# Gnd 0.01fF
C829 a_838_n225# Gnd 0.77fF
C830 p1 Gnd 13.73fF
C831 q6 Gnd 2.93fF
C832 qb1 Gnd 0.23fF
C833 a_17_n256# Gnd 0.16fF
C834 a1 Gnd 0.08fF
C835 a_55_n256# Gnd 0.23fF
C836 q1 Gnd 2.59fF
C837 a_110_n119# Gnd 0.01fF
C838 a_47_n115# Gnd 0.01fF
C839 a_281_n84# Gnd 0.01fF
C840 a_970_n61# Gnd 0.01fF
C841 c1 Gnd 0.08fF
C842 g0 Gnd 10.02fF
C843 qb5 Gnd 0.23fF
C844 a_17_n115# Gnd 0.16fF
C845 b0 Gnd 0.08fF
C846 g0_bar Gnd 9.56fF
C847 a_55_n115# Gnd 0.23fF
C848 a_874_36# Gnd 0.01fF
C849 qc0 Gnd 12.75fF
C850 a_841_36# Gnd 0.76fF
C851 a_243_2# Gnd 0.41fF
C852 a_112_19# Gnd 0.01fF
C853 a_49_23# Gnd 0.01fF
C854 gnd Gnd 44.44fF
C855 p0 Gnd 11.89fF
C856 qb0 Gnd 0.23fF
C857 rst Gnd 1.06fF
C858 a_19_23# Gnd 0.16fF
C859 clk Gnd 43.16fF
C860 a0 Gnd 0.08fF
C861 q5 Gnd 3.01fF
C862 a_57_23# Gnd 0.23fF
C863 q0 Gnd 2.47fF
C864 vdd Gnd 235.06fF

.tran 0.1n 700n

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))


run
plot v(clk)+14 v(rst)+12 v(c4)+8 v(c3)+6 v(c2)+4 v(c1)+2 v(cout)+10





.endc
.end
