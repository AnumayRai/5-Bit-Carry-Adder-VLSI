D Flip Flop
.include dff.cir
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

.param width_P= {20*lambda}
.param width_N= {10*lambda}
    
Vdd	vdd	gnd	'SUPPLY'
vclk clk gnd pulse 1.8 0 0ns 0ns 0ns 10ns 20ns
vin d gnd pwl 0 0 .2ns 1.8 13ns 1.8 14ns 0
vrst rst gnd PWL(0ns 0 30ns 0 31ns 1.8 700ns 1.8)

xdff_0 d clk rst q qb vdd gnd DFF
.tran 0.1n 200n

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))


run
plot v(clk)+8  v(rst)+6 v(d)+4 v(q)+2 

.endc
.end
