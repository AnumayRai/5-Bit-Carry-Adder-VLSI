magic
tech scmos
timestamp 1764648833
<< nwell >>
rect 6 40 163 101
rect 263 97 275 101
rect 230 57 326 97
rect 72 39 105 40
rect 230 20 254 57
rect 827 23 867 55
rect 4 -98 161 -37
rect 234 -97 274 -65
rect 332 -79 356 -42
rect 923 -74 963 -42
rect 70 -99 103 -98
rect 4 -239 161 -178
rect 263 -186 275 -182
rect 230 -226 326 -186
rect 70 -240 103 -239
rect 230 -263 254 -226
rect 824 -238 864 -206
rect 1010 -267 1050 -227
rect 818 -312 858 -272
rect 4 -381 161 -320
rect 234 -380 274 -348
rect 335 -367 359 -330
rect 70 -382 103 -381
rect 4 -568 161 -507
rect 263 -515 275 -511
rect 832 -512 872 -480
rect 230 -555 326 -515
rect 70 -569 103 -568
rect 230 -592 254 -555
rect 826 -586 866 -546
rect 1019 -606 1059 -558
rect 4 -710 161 -649
rect 234 -709 274 -677
rect 335 -693 359 -656
rect 826 -676 866 -628
rect 70 -711 103 -710
rect 834 -926 874 -894
rect 4 -1058 161 -997
rect 828 -1000 868 -960
rect 261 -1004 273 -1000
rect 228 -1044 324 -1004
rect 70 -1059 103 -1058
rect 228 -1081 252 -1044
rect 828 -1090 868 -1042
rect 1044 -1069 1084 -1013
rect 2 -1199 159 -1138
rect 232 -1198 272 -1166
rect 334 -1178 358 -1141
rect 829 -1185 869 -1129
rect 68 -1200 101 -1199
rect 833 -1421 873 -1389
rect 2 -1548 159 -1487
rect 260 -1494 272 -1490
rect 227 -1534 323 -1494
rect 827 -1495 867 -1455
rect 68 -1549 101 -1548
rect 227 -1571 251 -1534
rect 827 -1585 867 -1537
rect 1051 -1585 1091 -1521
rect 2 -1689 159 -1628
rect 231 -1688 271 -1656
rect 334 -1664 358 -1627
rect 828 -1680 868 -1624
rect 68 -1690 101 -1689
rect 824 -1792 864 -1728
rect 2 -2018 159 -1957
rect 68 -2019 101 -2018
<< ntransistor >>
rect 17 23 19 33
rect 47 23 49 33
rect 55 23 57 33
rect 110 19 112 29
rect 118 19 120 29
rect 150 22 152 32
rect 265 40 267 50
rect 288 34 290 44
rect 874 42 894 44
rect 874 34 894 36
rect 241 2 243 12
rect 970 -55 990 -53
rect 970 -63 990 -61
rect 281 -78 301 -76
rect 281 -86 301 -84
rect 15 -115 17 -105
rect 45 -115 47 -105
rect 53 -115 55 -105
rect 343 -97 345 -87
rect 108 -119 110 -109
rect 116 -119 118 -109
rect 148 -116 150 -106
rect 871 -219 891 -217
rect 871 -227 891 -225
rect 15 -256 17 -246
rect 45 -256 47 -246
rect 53 -256 55 -246
rect 108 -260 110 -250
rect 116 -260 118 -250
rect 148 -257 150 -247
rect 265 -243 267 -233
rect 288 -249 290 -239
rect 1057 -240 1087 -238
rect 1057 -248 1087 -246
rect 1057 -256 1087 -254
rect 241 -281 243 -271
rect 865 -285 895 -283
rect 865 -293 895 -291
rect 865 -301 895 -299
rect 281 -361 301 -359
rect 281 -369 301 -367
rect 15 -398 17 -388
rect 45 -398 47 -388
rect 53 -398 55 -388
rect 346 -385 348 -375
rect 108 -402 110 -392
rect 116 -402 118 -392
rect 148 -399 150 -389
rect 879 -493 899 -491
rect 879 -501 899 -499
rect 873 -559 903 -557
rect 15 -585 17 -575
rect 45 -585 47 -575
rect 53 -585 55 -575
rect 108 -589 110 -579
rect 116 -589 118 -579
rect 148 -586 150 -576
rect 265 -572 267 -562
rect 873 -567 903 -565
rect 288 -578 290 -568
rect 1066 -571 1106 -569
rect 873 -575 903 -573
rect 1066 -579 1106 -577
rect 1066 -587 1106 -585
rect 1066 -595 1106 -593
rect 241 -610 243 -600
rect 873 -641 913 -639
rect 873 -649 913 -647
rect 873 -657 913 -655
rect 873 -665 913 -663
rect 281 -690 301 -688
rect 281 -698 301 -696
rect 15 -727 17 -717
rect 45 -727 47 -717
rect 53 -727 55 -717
rect 346 -711 348 -701
rect 108 -731 110 -721
rect 116 -731 118 -721
rect 148 -728 150 -718
rect 881 -907 901 -905
rect 881 -915 901 -913
rect 875 -973 905 -971
rect 875 -981 905 -979
rect 875 -989 905 -987
rect 1091 -1026 1141 -1024
rect 1091 -1034 1141 -1032
rect 1091 -1042 1141 -1040
rect 15 -1075 17 -1065
rect 45 -1075 47 -1065
rect 53 -1075 55 -1065
rect 108 -1079 110 -1069
rect 116 -1079 118 -1069
rect 148 -1076 150 -1066
rect 263 -1061 265 -1051
rect 1091 -1050 1141 -1048
rect 875 -1055 915 -1053
rect 286 -1067 288 -1057
rect 1091 -1058 1141 -1056
rect 875 -1063 915 -1061
rect 875 -1071 915 -1069
rect 875 -1079 915 -1077
rect 239 -1099 241 -1089
rect 876 -1142 926 -1140
rect 876 -1150 926 -1148
rect 876 -1158 926 -1156
rect 876 -1166 926 -1164
rect 279 -1179 299 -1177
rect 279 -1187 299 -1185
rect 876 -1174 926 -1172
rect 13 -1216 15 -1206
rect 43 -1216 45 -1206
rect 51 -1216 53 -1206
rect 345 -1196 347 -1186
rect 106 -1220 108 -1210
rect 114 -1220 116 -1210
rect 146 -1217 148 -1207
rect 880 -1402 900 -1400
rect 880 -1410 900 -1408
rect 874 -1468 904 -1466
rect 874 -1476 904 -1474
rect 874 -1484 904 -1482
rect 1098 -1534 1158 -1532
rect 13 -1565 15 -1555
rect 43 -1565 45 -1555
rect 51 -1565 53 -1555
rect 106 -1569 108 -1559
rect 114 -1569 116 -1559
rect 146 -1566 148 -1556
rect 262 -1551 264 -1541
rect 1098 -1542 1158 -1540
rect 285 -1557 287 -1547
rect 874 -1550 914 -1548
rect 1098 -1550 1158 -1548
rect 874 -1558 914 -1556
rect 1098 -1558 1158 -1556
rect 874 -1566 914 -1564
rect 1098 -1566 1158 -1564
rect 874 -1574 914 -1572
rect 1098 -1574 1158 -1572
rect 238 -1589 240 -1579
rect 875 -1637 925 -1635
rect 875 -1645 925 -1643
rect 875 -1653 925 -1651
rect 278 -1669 298 -1667
rect 875 -1661 925 -1659
rect 875 -1669 925 -1667
rect 278 -1677 298 -1675
rect 345 -1682 347 -1672
rect 13 -1706 15 -1696
rect 43 -1706 45 -1696
rect 51 -1706 53 -1696
rect 106 -1710 108 -1700
rect 114 -1710 116 -1700
rect 146 -1707 148 -1697
rect 871 -1741 931 -1739
rect 871 -1749 931 -1747
rect 871 -1757 931 -1755
rect 871 -1765 931 -1763
rect 871 -1773 931 -1771
rect 871 -1781 931 -1779
rect 13 -2035 15 -2025
rect 43 -2035 45 -2025
rect 51 -2035 53 -2025
rect 106 -2039 108 -2029
rect 114 -2039 116 -2029
rect 146 -2036 148 -2026
<< ptransistor >>
rect 17 46 19 66
rect 25 46 27 66
rect 47 46 49 66
rect 55 46 57 66
rect 87 49 89 69
rect 110 62 112 82
rect 150 46 152 66
rect 265 63 267 83
rect 288 63 290 83
rect 241 26 243 46
rect 841 42 861 44
rect 841 34 861 36
rect 15 -92 17 -72
rect 23 -92 25 -72
rect 45 -92 47 -72
rect 53 -92 55 -72
rect 85 -89 87 -69
rect 108 -76 110 -56
rect 148 -92 150 -72
rect 343 -73 345 -53
rect 937 -55 957 -53
rect 937 -63 957 -61
rect 248 -78 268 -76
rect 248 -86 268 -84
rect 15 -233 17 -213
rect 23 -233 25 -213
rect 45 -233 47 -213
rect 53 -233 55 -213
rect 85 -230 87 -210
rect 108 -217 110 -197
rect 148 -233 150 -213
rect 265 -220 267 -200
rect 288 -220 290 -200
rect 838 -219 858 -217
rect 838 -227 858 -225
rect 241 -257 243 -237
rect 1024 -240 1044 -238
rect 1024 -248 1044 -246
rect 1024 -256 1044 -254
rect 832 -285 852 -283
rect 832 -293 852 -291
rect 832 -301 852 -299
rect 15 -375 17 -355
rect 23 -375 25 -355
rect 45 -375 47 -355
rect 53 -375 55 -355
rect 85 -372 87 -352
rect 108 -359 110 -339
rect 148 -375 150 -355
rect 248 -361 268 -359
rect 346 -361 348 -341
rect 248 -369 268 -367
rect 846 -493 866 -491
rect 846 -501 866 -499
rect 15 -562 17 -542
rect 23 -562 25 -542
rect 45 -562 47 -542
rect 53 -562 55 -542
rect 85 -559 87 -539
rect 108 -546 110 -526
rect 148 -562 150 -542
rect 265 -549 267 -529
rect 288 -549 290 -529
rect 840 -559 860 -557
rect 241 -586 243 -566
rect 840 -567 860 -565
rect 1033 -571 1053 -569
rect 840 -575 860 -573
rect 1033 -579 1053 -577
rect 1033 -587 1053 -585
rect 1033 -595 1053 -593
rect 840 -641 860 -639
rect 840 -649 860 -647
rect 840 -657 860 -655
rect 840 -665 860 -663
rect 15 -704 17 -684
rect 23 -704 25 -684
rect 45 -704 47 -684
rect 53 -704 55 -684
rect 85 -701 87 -681
rect 108 -688 110 -668
rect 148 -704 150 -684
rect 346 -687 348 -667
rect 248 -690 268 -688
rect 248 -698 268 -696
rect 848 -907 868 -905
rect 848 -915 868 -913
rect 842 -973 862 -971
rect 842 -981 862 -979
rect 842 -989 862 -987
rect 15 -1052 17 -1032
rect 23 -1052 25 -1032
rect 45 -1052 47 -1032
rect 53 -1052 55 -1032
rect 85 -1049 87 -1029
rect 108 -1036 110 -1016
rect 148 -1052 150 -1032
rect 263 -1038 265 -1018
rect 286 -1038 288 -1018
rect 1064 -1026 1078 -1024
rect 1064 -1034 1078 -1032
rect 1064 -1042 1078 -1040
rect 239 -1075 241 -1055
rect 1064 -1050 1078 -1048
rect 842 -1055 862 -1053
rect 1064 -1058 1078 -1056
rect 842 -1063 862 -1061
rect 842 -1071 862 -1069
rect 842 -1079 862 -1077
rect 849 -1142 863 -1140
rect 849 -1150 863 -1148
rect 13 -1193 15 -1173
rect 21 -1193 23 -1173
rect 43 -1193 45 -1173
rect 51 -1193 53 -1173
rect 83 -1190 85 -1170
rect 106 -1177 108 -1157
rect 345 -1172 347 -1152
rect 849 -1158 863 -1156
rect 849 -1166 863 -1164
rect 146 -1193 148 -1173
rect 246 -1179 266 -1177
rect 246 -1187 266 -1185
rect 849 -1174 863 -1172
rect 847 -1402 867 -1400
rect 847 -1410 867 -1408
rect 841 -1468 861 -1466
rect 841 -1476 861 -1474
rect 841 -1484 861 -1482
rect 13 -1542 15 -1522
rect 21 -1542 23 -1522
rect 43 -1542 45 -1522
rect 51 -1542 53 -1522
rect 83 -1539 85 -1519
rect 106 -1526 108 -1506
rect 146 -1542 148 -1522
rect 262 -1528 264 -1508
rect 285 -1528 287 -1508
rect 1065 -1534 1085 -1532
rect 238 -1565 240 -1545
rect 1065 -1542 1085 -1540
rect 841 -1550 861 -1548
rect 1065 -1550 1085 -1548
rect 841 -1558 861 -1556
rect 1065 -1558 1085 -1556
rect 841 -1566 861 -1564
rect 1065 -1566 1085 -1564
rect 841 -1574 861 -1572
rect 1065 -1574 1085 -1572
rect 848 -1637 862 -1635
rect 13 -1683 15 -1663
rect 21 -1683 23 -1663
rect 43 -1683 45 -1663
rect 51 -1683 53 -1663
rect 83 -1680 85 -1660
rect 106 -1667 108 -1647
rect 345 -1658 347 -1638
rect 848 -1645 862 -1643
rect 848 -1653 862 -1651
rect 146 -1683 148 -1663
rect 245 -1669 265 -1667
rect 848 -1661 862 -1659
rect 848 -1669 862 -1667
rect 245 -1677 265 -1675
rect 838 -1741 858 -1739
rect 838 -1749 858 -1747
rect 838 -1757 858 -1755
rect 838 -1765 858 -1763
rect 838 -1773 858 -1771
rect 838 -1781 858 -1779
rect 13 -2012 15 -1992
rect 21 -2012 23 -1992
rect 43 -2012 45 -1992
rect 51 -2012 53 -1992
rect 83 -2009 85 -1989
rect 106 -1996 108 -1976
rect 146 -2012 148 -1992
<< ndiffusion >>
rect 16 23 17 33
rect 19 23 20 33
rect 46 23 47 33
rect 49 23 50 33
rect 54 23 55 33
rect 57 23 58 33
rect 109 19 110 29
rect 112 19 113 29
rect 117 19 118 29
rect 120 19 121 29
rect 149 22 150 32
rect 152 22 153 32
rect 264 40 265 50
rect 267 40 268 50
rect 287 34 288 44
rect 290 34 291 44
rect 874 44 894 45
rect 874 41 894 42
rect 874 36 894 37
rect 874 33 894 34
rect 240 2 241 12
rect 243 2 244 12
rect 970 -53 990 -52
rect 970 -56 990 -55
rect 970 -61 990 -60
rect 970 -64 990 -63
rect 281 -76 301 -75
rect 281 -79 301 -78
rect 281 -84 301 -83
rect 281 -87 301 -86
rect 14 -115 15 -105
rect 17 -115 18 -105
rect 44 -115 45 -105
rect 47 -115 48 -105
rect 52 -115 53 -105
rect 55 -115 56 -105
rect 342 -97 343 -87
rect 345 -97 346 -87
rect 107 -119 108 -109
rect 110 -119 111 -109
rect 115 -119 116 -109
rect 118 -119 119 -109
rect 147 -116 148 -106
rect 150 -116 151 -106
rect 871 -217 891 -216
rect 871 -220 891 -219
rect 871 -225 891 -224
rect 871 -228 891 -227
rect 14 -256 15 -246
rect 17 -256 18 -246
rect 44 -256 45 -246
rect 47 -256 48 -246
rect 52 -256 53 -246
rect 55 -256 56 -246
rect 107 -260 108 -250
rect 110 -260 111 -250
rect 115 -260 116 -250
rect 118 -260 119 -250
rect 147 -257 148 -247
rect 150 -257 151 -247
rect 264 -243 265 -233
rect 267 -243 268 -233
rect 287 -249 288 -239
rect 290 -249 291 -239
rect 1057 -238 1087 -237
rect 1057 -241 1087 -240
rect 1057 -246 1087 -245
rect 1057 -249 1087 -248
rect 1057 -254 1087 -253
rect 1057 -257 1087 -256
rect 240 -281 241 -271
rect 243 -281 244 -271
rect 865 -283 895 -282
rect 865 -286 895 -285
rect 865 -291 895 -290
rect 865 -294 895 -293
rect 865 -299 895 -298
rect 865 -302 895 -301
rect 281 -359 301 -358
rect 281 -362 301 -361
rect 281 -367 301 -366
rect 281 -370 301 -369
rect 14 -398 15 -388
rect 17 -398 18 -388
rect 44 -398 45 -388
rect 47 -398 48 -388
rect 52 -398 53 -388
rect 55 -398 56 -388
rect 345 -385 346 -375
rect 348 -385 349 -375
rect 107 -402 108 -392
rect 110 -402 111 -392
rect 115 -402 116 -392
rect 118 -402 119 -392
rect 147 -399 148 -389
rect 150 -399 151 -389
rect 879 -491 899 -490
rect 879 -494 899 -493
rect 879 -499 899 -498
rect 879 -502 899 -501
rect 873 -557 903 -556
rect 14 -585 15 -575
rect 17 -585 18 -575
rect 44 -585 45 -575
rect 47 -585 48 -575
rect 52 -585 53 -575
rect 55 -585 56 -575
rect 107 -589 108 -579
rect 110 -589 111 -579
rect 115 -589 116 -579
rect 118 -589 119 -579
rect 147 -586 148 -576
rect 150 -586 151 -576
rect 264 -572 265 -562
rect 267 -572 268 -562
rect 873 -560 903 -559
rect 873 -565 903 -564
rect 287 -578 288 -568
rect 290 -578 291 -568
rect 873 -568 903 -567
rect 1066 -569 1106 -568
rect 873 -573 903 -572
rect 873 -576 903 -575
rect 1066 -572 1106 -571
rect 1066 -577 1106 -576
rect 1066 -580 1106 -579
rect 1066 -585 1106 -584
rect 1066 -588 1106 -587
rect 1066 -593 1106 -592
rect 1066 -596 1106 -595
rect 240 -610 241 -600
rect 243 -610 244 -600
rect 873 -639 913 -638
rect 873 -642 913 -641
rect 873 -647 913 -646
rect 873 -650 913 -649
rect 873 -655 913 -654
rect 873 -658 913 -657
rect 873 -663 913 -662
rect 873 -666 913 -665
rect 281 -688 301 -687
rect 281 -691 301 -690
rect 281 -696 301 -695
rect 281 -699 301 -698
rect 14 -727 15 -717
rect 17 -727 18 -717
rect 44 -727 45 -717
rect 47 -727 48 -717
rect 52 -727 53 -717
rect 55 -727 56 -717
rect 345 -711 346 -701
rect 348 -711 349 -701
rect 107 -731 108 -721
rect 110 -731 111 -721
rect 115 -731 116 -721
rect 118 -731 119 -721
rect 147 -728 148 -718
rect 150 -728 151 -718
rect 881 -905 901 -904
rect 881 -908 901 -907
rect 881 -913 901 -912
rect 881 -916 901 -915
rect 875 -971 905 -970
rect 875 -974 905 -973
rect 875 -979 905 -978
rect 875 -982 905 -981
rect 875 -987 905 -986
rect 875 -990 905 -989
rect 1091 -1024 1141 -1023
rect 1091 -1027 1141 -1026
rect 1091 -1032 1141 -1031
rect 1091 -1035 1141 -1034
rect 1091 -1040 1141 -1039
rect 14 -1075 15 -1065
rect 17 -1075 18 -1065
rect 44 -1075 45 -1065
rect 47 -1075 48 -1065
rect 52 -1075 53 -1065
rect 55 -1075 56 -1065
rect 107 -1079 108 -1069
rect 110 -1079 111 -1069
rect 115 -1079 116 -1069
rect 118 -1079 119 -1069
rect 147 -1076 148 -1066
rect 150 -1076 151 -1066
rect 262 -1061 263 -1051
rect 265 -1061 266 -1051
rect 1091 -1043 1141 -1042
rect 1091 -1048 1141 -1047
rect 875 -1053 915 -1052
rect 285 -1067 286 -1057
rect 288 -1067 289 -1057
rect 875 -1056 915 -1055
rect 1091 -1051 1141 -1050
rect 1091 -1056 1141 -1055
rect 875 -1061 915 -1060
rect 1091 -1059 1141 -1058
rect 875 -1064 915 -1063
rect 875 -1069 915 -1068
rect 875 -1072 915 -1071
rect 875 -1077 915 -1076
rect 875 -1080 915 -1079
rect 238 -1099 239 -1089
rect 241 -1099 242 -1089
rect 876 -1140 926 -1139
rect 876 -1143 926 -1142
rect 876 -1148 926 -1147
rect 876 -1151 926 -1150
rect 876 -1156 926 -1155
rect 876 -1159 926 -1158
rect 876 -1164 926 -1163
rect 876 -1167 926 -1166
rect 876 -1172 926 -1171
rect 279 -1177 299 -1176
rect 279 -1180 299 -1179
rect 279 -1185 299 -1184
rect 876 -1175 926 -1174
rect 279 -1188 299 -1187
rect 12 -1216 13 -1206
rect 15 -1216 16 -1206
rect 42 -1216 43 -1206
rect 45 -1216 46 -1206
rect 50 -1216 51 -1206
rect 53 -1216 54 -1206
rect 344 -1196 345 -1186
rect 347 -1196 348 -1186
rect 105 -1220 106 -1210
rect 108 -1220 109 -1210
rect 113 -1220 114 -1210
rect 116 -1220 117 -1210
rect 145 -1217 146 -1207
rect 148 -1217 149 -1207
rect 880 -1400 900 -1399
rect 880 -1403 900 -1402
rect 880 -1408 900 -1407
rect 880 -1411 900 -1410
rect 874 -1466 904 -1465
rect 874 -1469 904 -1468
rect 874 -1474 904 -1473
rect 874 -1477 904 -1476
rect 874 -1482 904 -1481
rect 874 -1485 904 -1484
rect 1098 -1532 1158 -1531
rect 12 -1565 13 -1555
rect 15 -1565 16 -1555
rect 42 -1565 43 -1555
rect 45 -1565 46 -1555
rect 50 -1565 51 -1555
rect 53 -1565 54 -1555
rect 105 -1569 106 -1559
rect 108 -1569 109 -1559
rect 113 -1569 114 -1559
rect 116 -1569 117 -1559
rect 145 -1566 146 -1556
rect 148 -1566 149 -1556
rect 261 -1551 262 -1541
rect 264 -1551 265 -1541
rect 1098 -1535 1158 -1534
rect 1098 -1540 1158 -1539
rect 284 -1557 285 -1547
rect 287 -1557 288 -1547
rect 874 -1548 914 -1547
rect 1098 -1543 1158 -1542
rect 1098 -1548 1158 -1547
rect 874 -1551 914 -1550
rect 874 -1556 914 -1555
rect 1098 -1551 1158 -1550
rect 1098 -1556 1158 -1555
rect 874 -1559 914 -1558
rect 874 -1564 914 -1563
rect 1098 -1559 1158 -1558
rect 1098 -1564 1158 -1563
rect 874 -1567 914 -1566
rect 874 -1572 914 -1571
rect 1098 -1567 1158 -1566
rect 1098 -1572 1158 -1571
rect 874 -1575 914 -1574
rect 1098 -1575 1158 -1574
rect 237 -1589 238 -1579
rect 240 -1589 241 -1579
rect 875 -1635 925 -1634
rect 875 -1638 925 -1637
rect 875 -1643 925 -1642
rect 875 -1646 925 -1645
rect 875 -1651 925 -1650
rect 278 -1667 298 -1666
rect 278 -1670 298 -1669
rect 875 -1654 925 -1653
rect 875 -1659 925 -1658
rect 875 -1662 925 -1661
rect 875 -1667 925 -1666
rect 278 -1675 298 -1674
rect 278 -1678 298 -1677
rect 344 -1682 345 -1672
rect 347 -1682 348 -1672
rect 875 -1670 925 -1669
rect 12 -1706 13 -1696
rect 15 -1706 16 -1696
rect 42 -1706 43 -1696
rect 45 -1706 46 -1696
rect 50 -1706 51 -1696
rect 53 -1706 54 -1696
rect 105 -1710 106 -1700
rect 108 -1710 109 -1700
rect 113 -1710 114 -1700
rect 116 -1710 117 -1700
rect 145 -1707 146 -1697
rect 148 -1707 149 -1697
rect 871 -1739 931 -1738
rect 871 -1742 931 -1741
rect 871 -1747 931 -1746
rect 871 -1750 931 -1749
rect 871 -1755 931 -1754
rect 871 -1758 931 -1757
rect 871 -1763 931 -1762
rect 871 -1766 931 -1765
rect 871 -1771 931 -1770
rect 871 -1774 931 -1773
rect 871 -1779 931 -1778
rect 871 -1782 931 -1781
rect 12 -2035 13 -2025
rect 15 -2035 16 -2025
rect 42 -2035 43 -2025
rect 45 -2035 46 -2025
rect 50 -2035 51 -2025
rect 53 -2035 54 -2025
rect 105 -2039 106 -2029
rect 108 -2039 109 -2029
rect 113 -2039 114 -2029
rect 116 -2039 117 -2029
rect 145 -2036 146 -2026
rect 148 -2036 149 -2026
<< pdiffusion >>
rect 16 46 17 66
rect 19 46 20 66
rect 24 46 25 66
rect 27 46 28 66
rect 46 46 47 66
rect 49 46 50 66
rect 54 46 55 66
rect 57 46 58 66
rect 86 49 87 69
rect 89 49 90 69
rect 109 62 110 82
rect 112 62 113 82
rect 149 46 150 66
rect 152 46 153 66
rect 264 63 265 83
rect 267 63 268 83
rect 287 63 288 83
rect 290 63 291 83
rect 240 26 241 46
rect 243 26 244 46
rect 841 44 861 45
rect 841 41 861 42
rect 841 36 861 37
rect 841 33 861 34
rect 14 -92 15 -72
rect 17 -92 18 -72
rect 22 -92 23 -72
rect 25 -92 26 -72
rect 44 -92 45 -72
rect 47 -92 48 -72
rect 52 -92 53 -72
rect 55 -92 56 -72
rect 84 -89 85 -69
rect 87 -89 88 -69
rect 107 -76 108 -56
rect 110 -76 111 -56
rect 147 -92 148 -72
rect 150 -92 151 -72
rect 248 -76 268 -75
rect 342 -73 343 -53
rect 345 -73 346 -53
rect 937 -53 957 -52
rect 937 -56 957 -55
rect 937 -61 957 -60
rect 937 -64 957 -63
rect 248 -79 268 -78
rect 248 -84 268 -83
rect 248 -87 268 -86
rect 14 -233 15 -213
rect 17 -233 18 -213
rect 22 -233 23 -213
rect 25 -233 26 -213
rect 44 -233 45 -213
rect 47 -233 48 -213
rect 52 -233 53 -213
rect 55 -233 56 -213
rect 84 -230 85 -210
rect 87 -230 88 -210
rect 107 -217 108 -197
rect 110 -217 111 -197
rect 147 -233 148 -213
rect 150 -233 151 -213
rect 264 -220 265 -200
rect 267 -220 268 -200
rect 287 -220 288 -200
rect 290 -220 291 -200
rect 838 -217 858 -216
rect 838 -220 858 -219
rect 838 -225 858 -224
rect 838 -228 858 -227
rect 240 -257 241 -237
rect 243 -257 244 -237
rect 1024 -238 1044 -237
rect 1024 -241 1044 -240
rect 1024 -246 1044 -245
rect 1024 -249 1044 -248
rect 1024 -254 1044 -253
rect 1024 -257 1044 -256
rect 832 -283 852 -282
rect 832 -286 852 -285
rect 832 -291 852 -290
rect 832 -294 852 -293
rect 832 -299 852 -298
rect 832 -302 852 -301
rect 14 -375 15 -355
rect 17 -375 18 -355
rect 22 -375 23 -355
rect 25 -375 26 -355
rect 44 -375 45 -355
rect 47 -375 48 -355
rect 52 -375 53 -355
rect 55 -375 56 -355
rect 84 -372 85 -352
rect 87 -372 88 -352
rect 107 -359 108 -339
rect 110 -359 111 -339
rect 147 -375 148 -355
rect 150 -375 151 -355
rect 248 -359 268 -358
rect 345 -361 346 -341
rect 348 -361 349 -341
rect 248 -362 268 -361
rect 248 -367 268 -366
rect 248 -370 268 -369
rect 846 -491 866 -490
rect 846 -494 866 -493
rect 846 -499 866 -498
rect 846 -502 866 -501
rect 14 -562 15 -542
rect 17 -562 18 -542
rect 22 -562 23 -542
rect 25 -562 26 -542
rect 44 -562 45 -542
rect 47 -562 48 -542
rect 52 -562 53 -542
rect 55 -562 56 -542
rect 84 -559 85 -539
rect 87 -559 88 -539
rect 107 -546 108 -526
rect 110 -546 111 -526
rect 147 -562 148 -542
rect 150 -562 151 -542
rect 264 -549 265 -529
rect 267 -549 268 -529
rect 287 -549 288 -529
rect 290 -549 291 -529
rect 840 -557 860 -556
rect 840 -560 860 -559
rect 240 -586 241 -566
rect 243 -586 244 -566
rect 840 -565 860 -564
rect 840 -568 860 -567
rect 840 -573 860 -572
rect 1033 -569 1053 -568
rect 1033 -572 1053 -571
rect 840 -576 860 -575
rect 1033 -577 1053 -576
rect 1033 -580 1053 -579
rect 1033 -585 1053 -584
rect 1033 -588 1053 -587
rect 1033 -593 1053 -592
rect 1033 -596 1053 -595
rect 840 -639 860 -638
rect 840 -642 860 -641
rect 840 -647 860 -646
rect 840 -650 860 -649
rect 840 -655 860 -654
rect 840 -658 860 -657
rect 840 -663 860 -662
rect 840 -666 860 -665
rect 14 -704 15 -684
rect 17 -704 18 -684
rect 22 -704 23 -684
rect 25 -704 26 -684
rect 44 -704 45 -684
rect 47 -704 48 -684
rect 52 -704 53 -684
rect 55 -704 56 -684
rect 84 -701 85 -681
rect 87 -701 88 -681
rect 107 -688 108 -668
rect 110 -688 111 -668
rect 147 -704 148 -684
rect 150 -704 151 -684
rect 248 -688 268 -687
rect 345 -687 346 -667
rect 348 -687 349 -667
rect 248 -691 268 -690
rect 248 -696 268 -695
rect 248 -699 268 -698
rect 848 -905 868 -904
rect 848 -908 868 -907
rect 848 -913 868 -912
rect 848 -916 868 -915
rect 842 -971 862 -970
rect 842 -974 862 -973
rect 842 -979 862 -978
rect 842 -982 862 -981
rect 842 -987 862 -986
rect 842 -990 862 -989
rect 14 -1052 15 -1032
rect 17 -1052 18 -1032
rect 22 -1052 23 -1032
rect 25 -1052 26 -1032
rect 44 -1052 45 -1032
rect 47 -1052 48 -1032
rect 52 -1052 53 -1032
rect 55 -1052 56 -1032
rect 84 -1049 85 -1029
rect 87 -1049 88 -1029
rect 107 -1036 108 -1016
rect 110 -1036 111 -1016
rect 147 -1052 148 -1032
rect 150 -1052 151 -1032
rect 262 -1038 263 -1018
rect 265 -1038 266 -1018
rect 285 -1038 286 -1018
rect 288 -1038 289 -1018
rect 1064 -1024 1078 -1023
rect 1064 -1027 1078 -1026
rect 1064 -1032 1078 -1031
rect 1064 -1035 1078 -1034
rect 1064 -1040 1078 -1039
rect 1064 -1043 1078 -1042
rect 238 -1075 239 -1055
rect 241 -1075 242 -1055
rect 842 -1053 862 -1052
rect 1064 -1048 1078 -1047
rect 1064 -1051 1078 -1050
rect 842 -1056 862 -1055
rect 842 -1061 862 -1060
rect 1064 -1056 1078 -1055
rect 1064 -1059 1078 -1058
rect 842 -1064 862 -1063
rect 842 -1069 862 -1068
rect 842 -1072 862 -1071
rect 842 -1077 862 -1076
rect 842 -1080 862 -1079
rect 849 -1140 863 -1139
rect 849 -1143 863 -1142
rect 849 -1148 863 -1147
rect 849 -1151 863 -1150
rect 12 -1193 13 -1173
rect 15 -1193 16 -1173
rect 20 -1193 21 -1173
rect 23 -1193 24 -1173
rect 42 -1193 43 -1173
rect 45 -1193 46 -1173
rect 50 -1193 51 -1173
rect 53 -1193 54 -1173
rect 82 -1190 83 -1170
rect 85 -1190 86 -1170
rect 105 -1177 106 -1157
rect 108 -1177 109 -1157
rect 344 -1172 345 -1152
rect 347 -1172 348 -1152
rect 849 -1156 863 -1155
rect 849 -1159 863 -1158
rect 849 -1164 863 -1163
rect 849 -1167 863 -1166
rect 849 -1172 863 -1171
rect 145 -1193 146 -1173
rect 148 -1193 149 -1173
rect 246 -1177 266 -1176
rect 246 -1180 266 -1179
rect 246 -1185 266 -1184
rect 849 -1175 863 -1174
rect 246 -1188 266 -1187
rect 847 -1400 867 -1399
rect 847 -1403 867 -1402
rect 847 -1408 867 -1407
rect 847 -1411 867 -1410
rect 841 -1466 861 -1465
rect 841 -1469 861 -1468
rect 841 -1474 861 -1473
rect 841 -1477 861 -1476
rect 841 -1482 861 -1481
rect 841 -1485 861 -1484
rect 12 -1542 13 -1522
rect 15 -1542 16 -1522
rect 20 -1542 21 -1522
rect 23 -1542 24 -1522
rect 42 -1542 43 -1522
rect 45 -1542 46 -1522
rect 50 -1542 51 -1522
rect 53 -1542 54 -1522
rect 82 -1539 83 -1519
rect 85 -1539 86 -1519
rect 105 -1526 106 -1506
rect 108 -1526 109 -1506
rect 145 -1542 146 -1522
rect 148 -1542 149 -1522
rect 261 -1528 262 -1508
rect 264 -1528 265 -1508
rect 284 -1528 285 -1508
rect 287 -1528 288 -1508
rect 1065 -1532 1085 -1531
rect 1065 -1535 1085 -1534
rect 237 -1565 238 -1545
rect 240 -1565 241 -1545
rect 1065 -1540 1085 -1539
rect 1065 -1543 1085 -1542
rect 841 -1548 861 -1547
rect 1065 -1548 1085 -1547
rect 841 -1551 861 -1550
rect 841 -1556 861 -1555
rect 1065 -1551 1085 -1550
rect 1065 -1556 1085 -1555
rect 841 -1559 861 -1558
rect 841 -1564 861 -1563
rect 1065 -1559 1085 -1558
rect 1065 -1564 1085 -1563
rect 841 -1567 861 -1566
rect 841 -1572 861 -1571
rect 1065 -1567 1085 -1566
rect 1065 -1572 1085 -1571
rect 841 -1575 861 -1574
rect 1065 -1575 1085 -1574
rect 848 -1635 862 -1634
rect 848 -1638 862 -1637
rect 12 -1683 13 -1663
rect 15 -1683 16 -1663
rect 20 -1683 21 -1663
rect 23 -1683 24 -1663
rect 42 -1683 43 -1663
rect 45 -1683 46 -1663
rect 50 -1683 51 -1663
rect 53 -1683 54 -1663
rect 82 -1680 83 -1660
rect 85 -1680 86 -1660
rect 105 -1667 106 -1647
rect 108 -1667 109 -1647
rect 344 -1658 345 -1638
rect 347 -1658 348 -1638
rect 848 -1643 862 -1642
rect 848 -1646 862 -1645
rect 848 -1651 862 -1650
rect 848 -1654 862 -1653
rect 145 -1683 146 -1663
rect 148 -1683 149 -1663
rect 245 -1667 265 -1666
rect 245 -1670 265 -1669
rect 245 -1675 265 -1674
rect 848 -1659 862 -1658
rect 848 -1662 862 -1661
rect 848 -1667 862 -1666
rect 848 -1670 862 -1669
rect 245 -1678 265 -1677
rect 838 -1739 858 -1738
rect 838 -1742 858 -1741
rect 838 -1747 858 -1746
rect 838 -1750 858 -1749
rect 838 -1755 858 -1754
rect 838 -1758 858 -1757
rect 838 -1763 858 -1762
rect 838 -1766 858 -1765
rect 838 -1771 858 -1770
rect 838 -1774 858 -1773
rect 838 -1779 858 -1778
rect 838 -1782 858 -1781
rect 12 -2012 13 -1992
rect 15 -2012 16 -1992
rect 20 -2012 21 -1992
rect 23 -2012 24 -1992
rect 42 -2012 43 -1992
rect 45 -2012 46 -1992
rect 50 -2012 51 -1992
rect 53 -2012 54 -1992
rect 82 -2009 83 -1989
rect 85 -2009 86 -1989
rect 105 -1996 106 -1976
rect 108 -1996 109 -1976
rect 145 -2012 146 -1992
rect 148 -2012 149 -1992
<< ndcontact >>
rect 12 23 16 33
rect 20 23 32 33
rect 42 23 46 33
rect 50 23 54 33
rect 58 23 62 33
rect 105 19 109 29
rect 113 19 117 29
rect 121 19 125 29
rect 145 22 149 32
rect 153 22 157 32
rect 260 40 264 50
rect 268 40 272 50
rect 283 34 287 44
rect 291 34 295 44
rect 874 45 894 49
rect 874 37 894 41
rect 874 29 894 33
rect 236 2 240 12
rect 244 2 248 12
rect 281 -75 301 -71
rect 970 -52 990 -48
rect 970 -60 990 -56
rect 970 -68 990 -64
rect 281 -83 301 -79
rect 281 -91 301 -87
rect 10 -115 14 -105
rect 18 -115 30 -105
rect 40 -115 44 -105
rect 48 -115 52 -105
rect 56 -115 60 -105
rect 338 -97 342 -87
rect 346 -97 350 -87
rect 103 -119 107 -109
rect 111 -119 115 -109
rect 119 -119 123 -109
rect 143 -116 147 -106
rect 151 -116 155 -106
rect 871 -216 891 -212
rect 871 -224 891 -220
rect 871 -232 891 -228
rect 10 -256 14 -246
rect 18 -256 30 -246
rect 40 -256 44 -246
rect 48 -256 52 -246
rect 56 -256 60 -246
rect 103 -260 107 -250
rect 111 -260 115 -250
rect 119 -260 123 -250
rect 143 -257 147 -247
rect 151 -257 155 -247
rect 260 -243 264 -233
rect 268 -243 272 -233
rect 283 -249 287 -239
rect 291 -249 295 -239
rect 1057 -237 1087 -233
rect 1057 -245 1087 -241
rect 1057 -253 1087 -249
rect 1057 -261 1087 -257
rect 236 -281 240 -271
rect 244 -281 248 -271
rect 865 -282 895 -278
rect 865 -290 895 -286
rect 865 -298 895 -294
rect 865 -306 895 -302
rect 281 -358 301 -354
rect 281 -366 301 -362
rect 281 -374 301 -370
rect 10 -398 14 -388
rect 18 -398 30 -388
rect 40 -398 44 -388
rect 48 -398 52 -388
rect 56 -398 60 -388
rect 341 -385 345 -375
rect 349 -385 353 -375
rect 103 -402 107 -392
rect 111 -402 115 -392
rect 119 -402 123 -392
rect 143 -399 147 -389
rect 151 -399 155 -389
rect 879 -490 899 -486
rect 879 -498 899 -494
rect 879 -506 899 -502
rect 873 -556 903 -552
rect 10 -585 14 -575
rect 18 -585 30 -575
rect 40 -585 44 -575
rect 48 -585 52 -575
rect 56 -585 60 -575
rect 103 -589 107 -579
rect 111 -589 115 -579
rect 119 -589 123 -579
rect 143 -586 147 -576
rect 151 -586 155 -576
rect 260 -572 264 -562
rect 268 -572 272 -562
rect 873 -564 903 -560
rect 283 -578 287 -568
rect 291 -578 295 -568
rect 873 -572 903 -568
rect 1066 -568 1106 -564
rect 873 -580 903 -576
rect 1066 -576 1106 -572
rect 1066 -584 1106 -580
rect 1066 -592 1106 -588
rect 1066 -600 1106 -596
rect 236 -610 240 -600
rect 244 -610 248 -600
rect 873 -638 913 -634
rect 873 -646 913 -642
rect 873 -654 913 -650
rect 873 -662 913 -658
rect 281 -687 301 -683
rect 873 -670 913 -666
rect 281 -695 301 -691
rect 281 -703 301 -699
rect 10 -727 14 -717
rect 18 -727 30 -717
rect 40 -727 44 -717
rect 48 -727 52 -717
rect 56 -727 60 -717
rect 341 -711 345 -701
rect 349 -711 353 -701
rect 103 -731 107 -721
rect 111 -731 115 -721
rect 119 -731 123 -721
rect 143 -728 147 -718
rect 151 -728 155 -718
rect 881 -904 901 -900
rect 881 -912 901 -908
rect 881 -920 901 -916
rect 875 -970 905 -966
rect 875 -978 905 -974
rect 875 -986 905 -982
rect 875 -994 905 -990
rect 1091 -1023 1141 -1019
rect 1091 -1031 1141 -1027
rect 1091 -1039 1141 -1035
rect 10 -1075 14 -1065
rect 18 -1075 30 -1065
rect 40 -1075 44 -1065
rect 48 -1075 52 -1065
rect 56 -1075 60 -1065
rect 103 -1079 107 -1069
rect 111 -1079 115 -1069
rect 119 -1079 123 -1069
rect 143 -1076 147 -1066
rect 151 -1076 155 -1066
rect 258 -1061 262 -1051
rect 266 -1061 270 -1051
rect 875 -1052 915 -1048
rect 1091 -1047 1141 -1043
rect 281 -1067 285 -1057
rect 289 -1067 293 -1057
rect 875 -1060 915 -1056
rect 1091 -1055 1141 -1051
rect 1091 -1063 1141 -1059
rect 875 -1068 915 -1064
rect 875 -1076 915 -1072
rect 875 -1084 915 -1080
rect 234 -1099 238 -1089
rect 242 -1099 246 -1089
rect 876 -1139 926 -1135
rect 876 -1147 926 -1143
rect 876 -1155 926 -1151
rect 876 -1163 926 -1159
rect 876 -1171 926 -1167
rect 279 -1176 299 -1172
rect 279 -1184 299 -1180
rect 876 -1179 926 -1175
rect 279 -1192 299 -1188
rect 8 -1216 12 -1206
rect 16 -1216 28 -1206
rect 38 -1216 42 -1206
rect 46 -1216 50 -1206
rect 54 -1216 58 -1206
rect 340 -1196 344 -1186
rect 348 -1196 352 -1186
rect 101 -1220 105 -1210
rect 109 -1220 113 -1210
rect 117 -1220 121 -1210
rect 141 -1217 145 -1207
rect 149 -1217 153 -1207
rect 880 -1399 900 -1395
rect 880 -1407 900 -1403
rect 880 -1415 900 -1411
rect 874 -1465 904 -1461
rect 874 -1473 904 -1469
rect 874 -1481 904 -1477
rect 874 -1489 904 -1485
rect 1098 -1531 1158 -1527
rect 8 -1565 12 -1555
rect 16 -1565 28 -1555
rect 38 -1565 42 -1555
rect 46 -1565 50 -1555
rect 54 -1565 58 -1555
rect 101 -1569 105 -1559
rect 109 -1569 113 -1559
rect 117 -1569 121 -1559
rect 141 -1566 145 -1556
rect 149 -1566 153 -1556
rect 257 -1551 261 -1541
rect 265 -1551 269 -1541
rect 1098 -1539 1158 -1535
rect 280 -1557 284 -1547
rect 288 -1557 292 -1547
rect 874 -1547 914 -1543
rect 1098 -1547 1158 -1543
rect 874 -1555 914 -1551
rect 1098 -1555 1158 -1551
rect 874 -1563 914 -1559
rect 1098 -1563 1158 -1559
rect 874 -1571 914 -1567
rect 1098 -1571 1158 -1567
rect 874 -1579 914 -1575
rect 1098 -1579 1158 -1575
rect 233 -1589 237 -1579
rect 241 -1589 245 -1579
rect 875 -1634 925 -1630
rect 875 -1642 925 -1638
rect 875 -1650 925 -1646
rect 278 -1666 298 -1662
rect 278 -1674 298 -1670
rect 875 -1658 925 -1654
rect 875 -1666 925 -1662
rect 278 -1682 298 -1678
rect 340 -1682 344 -1672
rect 348 -1682 352 -1672
rect 875 -1674 925 -1670
rect 8 -1706 12 -1696
rect 16 -1706 28 -1696
rect 38 -1706 42 -1696
rect 46 -1706 50 -1696
rect 54 -1706 58 -1696
rect 101 -1710 105 -1700
rect 109 -1710 113 -1700
rect 117 -1710 121 -1700
rect 141 -1707 145 -1697
rect 149 -1707 153 -1697
rect 871 -1738 931 -1734
rect 871 -1746 931 -1742
rect 871 -1754 931 -1750
rect 871 -1762 931 -1758
rect 871 -1770 931 -1766
rect 871 -1778 931 -1774
rect 871 -1786 931 -1782
rect 8 -2035 12 -2025
rect 16 -2035 28 -2025
rect 38 -2035 42 -2025
rect 46 -2035 50 -2025
rect 54 -2035 58 -2025
rect 101 -2039 105 -2029
rect 109 -2039 113 -2029
rect 117 -2039 121 -2029
rect 141 -2036 145 -2026
rect 149 -2036 153 -2026
<< pdcontact >>
rect 12 46 16 66
rect 20 46 24 66
rect 28 46 32 66
rect 42 46 46 66
rect 50 46 54 66
rect 58 46 62 66
rect 82 49 86 69
rect 90 49 94 69
rect 105 62 109 82
rect 113 62 125 82
rect 145 46 149 66
rect 153 46 157 66
rect 260 63 264 83
rect 268 63 272 83
rect 283 63 287 83
rect 291 63 295 83
rect 236 26 240 46
rect 244 26 248 46
rect 841 45 861 49
rect 841 37 861 41
rect 841 29 861 33
rect 10 -92 14 -72
rect 18 -92 22 -72
rect 26 -92 30 -72
rect 40 -92 44 -72
rect 48 -92 52 -72
rect 56 -92 60 -72
rect 80 -89 84 -69
rect 88 -89 92 -69
rect 103 -76 107 -56
rect 111 -76 123 -56
rect 143 -92 147 -72
rect 151 -92 155 -72
rect 248 -75 268 -71
rect 338 -73 342 -53
rect 346 -73 350 -53
rect 937 -52 957 -48
rect 937 -60 957 -56
rect 937 -68 957 -64
rect 248 -83 268 -79
rect 248 -91 268 -87
rect 10 -233 14 -213
rect 18 -233 22 -213
rect 26 -233 30 -213
rect 40 -233 44 -213
rect 48 -233 52 -213
rect 56 -233 60 -213
rect 80 -230 84 -210
rect 88 -230 92 -210
rect 103 -217 107 -197
rect 111 -217 123 -197
rect 143 -233 147 -213
rect 151 -233 155 -213
rect 260 -220 264 -200
rect 268 -220 272 -200
rect 283 -220 287 -200
rect 291 -220 295 -200
rect 838 -216 858 -212
rect 838 -224 858 -220
rect 838 -232 858 -228
rect 236 -257 240 -237
rect 244 -257 248 -237
rect 1024 -237 1044 -233
rect 1024 -245 1044 -241
rect 1024 -253 1044 -249
rect 1024 -261 1044 -257
rect 832 -282 852 -278
rect 832 -290 852 -286
rect 832 -298 852 -294
rect 832 -306 852 -302
rect 10 -375 14 -355
rect 18 -375 22 -355
rect 26 -375 30 -355
rect 40 -375 44 -355
rect 48 -375 52 -355
rect 56 -375 60 -355
rect 80 -372 84 -352
rect 88 -372 92 -352
rect 103 -359 107 -339
rect 111 -359 123 -339
rect 143 -375 147 -355
rect 151 -375 155 -355
rect 248 -358 268 -354
rect 341 -361 345 -341
rect 349 -361 353 -341
rect 248 -366 268 -362
rect 248 -374 268 -370
rect 846 -490 866 -486
rect 846 -498 866 -494
rect 846 -506 866 -502
rect 10 -562 14 -542
rect 18 -562 22 -542
rect 26 -562 30 -542
rect 40 -562 44 -542
rect 48 -562 52 -542
rect 56 -562 60 -542
rect 80 -559 84 -539
rect 88 -559 92 -539
rect 103 -546 107 -526
rect 111 -546 123 -526
rect 143 -562 147 -542
rect 151 -562 155 -542
rect 260 -549 264 -529
rect 268 -549 272 -529
rect 283 -549 287 -529
rect 291 -549 295 -529
rect 840 -556 860 -552
rect 236 -586 240 -566
rect 244 -586 248 -566
rect 840 -564 860 -560
rect 840 -572 860 -568
rect 1033 -568 1053 -564
rect 840 -580 860 -576
rect 1033 -576 1053 -572
rect 1033 -584 1053 -580
rect 1033 -592 1053 -588
rect 1033 -600 1053 -596
rect 840 -638 860 -634
rect 840 -646 860 -642
rect 840 -654 860 -650
rect 840 -662 860 -658
rect 10 -704 14 -684
rect 18 -704 22 -684
rect 26 -704 30 -684
rect 40 -704 44 -684
rect 48 -704 52 -684
rect 56 -704 60 -684
rect 80 -701 84 -681
rect 88 -701 92 -681
rect 103 -688 107 -668
rect 111 -688 123 -668
rect 143 -704 147 -684
rect 151 -704 155 -684
rect 248 -687 268 -683
rect 341 -687 345 -667
rect 349 -687 353 -667
rect 840 -670 860 -666
rect 248 -695 268 -691
rect 248 -703 268 -699
rect 848 -904 868 -900
rect 848 -912 868 -908
rect 848 -920 868 -916
rect 842 -970 862 -966
rect 842 -978 862 -974
rect 842 -986 862 -982
rect 842 -994 862 -990
rect 10 -1052 14 -1032
rect 18 -1052 22 -1032
rect 26 -1052 30 -1032
rect 40 -1052 44 -1032
rect 48 -1052 52 -1032
rect 56 -1052 60 -1032
rect 80 -1049 84 -1029
rect 88 -1049 92 -1029
rect 103 -1036 107 -1016
rect 111 -1036 123 -1016
rect 143 -1052 147 -1032
rect 151 -1052 155 -1032
rect 258 -1038 262 -1018
rect 266 -1038 270 -1018
rect 281 -1038 285 -1018
rect 289 -1038 293 -1018
rect 1064 -1023 1078 -1019
rect 1064 -1031 1078 -1027
rect 1064 -1039 1078 -1035
rect 1064 -1047 1078 -1043
rect 234 -1075 238 -1055
rect 242 -1075 246 -1055
rect 842 -1052 862 -1048
rect 1064 -1055 1078 -1051
rect 842 -1060 862 -1056
rect 1064 -1063 1078 -1059
rect 842 -1068 862 -1064
rect 842 -1076 862 -1072
rect 842 -1084 862 -1080
rect 849 -1139 863 -1135
rect 849 -1147 863 -1143
rect 8 -1193 12 -1173
rect 16 -1193 20 -1173
rect 24 -1193 28 -1173
rect 38 -1193 42 -1173
rect 46 -1193 50 -1173
rect 54 -1193 58 -1173
rect 78 -1190 82 -1170
rect 86 -1190 90 -1170
rect 101 -1177 105 -1157
rect 109 -1177 121 -1157
rect 340 -1172 344 -1152
rect 348 -1172 352 -1152
rect 849 -1155 863 -1151
rect 849 -1163 863 -1159
rect 849 -1171 863 -1167
rect 141 -1193 145 -1173
rect 149 -1193 153 -1173
rect 246 -1176 266 -1172
rect 246 -1184 266 -1180
rect 849 -1179 863 -1175
rect 246 -1192 266 -1188
rect 847 -1399 867 -1395
rect 847 -1407 867 -1403
rect 847 -1415 867 -1411
rect 841 -1465 861 -1461
rect 841 -1473 861 -1469
rect 841 -1481 861 -1477
rect 841 -1489 861 -1485
rect 8 -1542 12 -1522
rect 16 -1542 20 -1522
rect 24 -1542 28 -1522
rect 38 -1542 42 -1522
rect 46 -1542 50 -1522
rect 54 -1542 58 -1522
rect 78 -1539 82 -1519
rect 86 -1539 90 -1519
rect 101 -1526 105 -1506
rect 109 -1526 121 -1506
rect 141 -1542 145 -1522
rect 149 -1542 153 -1522
rect 257 -1528 261 -1508
rect 265 -1528 269 -1508
rect 280 -1528 284 -1508
rect 288 -1528 292 -1508
rect 1065 -1531 1085 -1527
rect 233 -1565 237 -1545
rect 241 -1565 245 -1545
rect 1065 -1539 1085 -1535
rect 841 -1547 861 -1543
rect 1065 -1547 1085 -1543
rect 841 -1555 861 -1551
rect 1065 -1555 1085 -1551
rect 841 -1563 861 -1559
rect 1065 -1563 1085 -1559
rect 841 -1571 861 -1567
rect 1065 -1571 1085 -1567
rect 841 -1579 861 -1575
rect 1065 -1579 1085 -1575
rect 848 -1634 862 -1630
rect 8 -1683 12 -1663
rect 16 -1683 20 -1663
rect 24 -1683 28 -1663
rect 38 -1683 42 -1663
rect 46 -1683 50 -1663
rect 54 -1683 58 -1663
rect 78 -1680 82 -1660
rect 86 -1680 90 -1660
rect 101 -1667 105 -1647
rect 109 -1667 121 -1647
rect 340 -1658 344 -1638
rect 348 -1658 352 -1638
rect 848 -1642 862 -1638
rect 848 -1650 862 -1646
rect 848 -1658 862 -1654
rect 141 -1683 145 -1663
rect 149 -1683 153 -1663
rect 245 -1666 265 -1662
rect 245 -1674 265 -1670
rect 848 -1666 862 -1662
rect 245 -1682 265 -1678
rect 848 -1674 862 -1670
rect 838 -1738 858 -1734
rect 838 -1746 858 -1742
rect 838 -1754 858 -1750
rect 838 -1762 858 -1758
rect 838 -1770 858 -1766
rect 838 -1778 858 -1774
rect 838 -1786 858 -1782
rect 8 -2012 12 -1992
rect 16 -2012 20 -1992
rect 24 -2012 28 -1992
rect 38 -2012 42 -1992
rect 46 -2012 50 -1992
rect 54 -2012 58 -1992
rect 78 -2009 82 -1989
rect 86 -2009 90 -1989
rect 101 -1996 105 -1976
rect 109 -1996 121 -1976
rect 141 -2012 145 -1992
rect 149 -2012 153 -1992
<< psubstratepcontact >>
rect 0 0 4 5
rect 236 -6 240 -2
rect 305 -91 309 -87
rect 338 -105 342 -101
rect -2 -138 2 -133
rect -2 -279 2 -274
rect 236 -289 240 -285
rect 305 -374 309 -370
rect 341 -393 345 -389
rect -2 -421 2 -416
rect -2 -608 2 -603
rect 236 -618 240 -614
rect 305 -703 309 -699
rect 341 -719 345 -715
rect -2 -750 2 -745
rect -2 -1098 2 -1093
rect 234 -1107 238 -1103
rect 303 -1192 307 -1188
rect 340 -1204 344 -1200
rect -4 -1239 0 -1234
rect -4 -1588 0 -1583
rect 233 -1597 237 -1593
rect 302 -1682 306 -1678
rect 340 -1690 344 -1686
rect -4 -1729 0 -1724
rect -4 -2058 0 -2053
<< nsubstratencontact >>
rect 155 90 159 94
rect 236 50 240 54
rect 832 29 836 33
rect 153 -48 157 -44
rect 338 -49 342 -45
rect 928 -68 932 -64
rect 239 -91 243 -87
rect 153 -189 157 -185
rect 236 -233 240 -229
rect 829 -232 833 -228
rect 1015 -261 1019 -257
rect 823 -306 827 -302
rect 153 -331 157 -327
rect 341 -337 345 -333
rect 239 -374 243 -370
rect 837 -506 841 -502
rect 153 -518 157 -514
rect 236 -562 240 -558
rect 831 -580 835 -576
rect 1024 -600 1028 -596
rect 153 -660 157 -656
rect 341 -663 345 -659
rect 831 -670 835 -666
rect 239 -703 243 -699
rect 839 -920 843 -916
rect 833 -994 837 -990
rect 153 -1008 157 -1004
rect 234 -1051 238 -1047
rect 1051 -1063 1055 -1059
rect 833 -1084 837 -1080
rect 151 -1149 155 -1145
rect 340 -1148 344 -1144
rect 836 -1179 840 -1175
rect 237 -1192 241 -1188
rect 838 -1415 842 -1411
rect 832 -1489 836 -1485
rect 151 -1498 155 -1494
rect 233 -1541 237 -1537
rect 832 -1579 836 -1575
rect 1056 -1579 1060 -1575
rect 340 -1634 344 -1630
rect 151 -1639 155 -1635
rect 236 -1682 240 -1678
rect 835 -1674 839 -1670
rect 829 -1786 833 -1782
rect 151 -1968 155 -1964
<< polysilicon >>
rect 110 82 112 86
rect 265 83 267 96
rect 288 83 290 87
rect 17 66 19 70
rect 25 66 27 70
rect 47 66 49 70
rect 55 66 57 70
rect 87 69 89 73
rect 150 66 152 70
rect 17 33 19 46
rect 25 42 27 46
rect 47 33 49 46
rect 55 33 57 46
rect 87 45 89 49
rect 110 43 112 62
rect 265 50 267 63
rect 288 59 290 63
rect 241 46 243 49
rect 110 29 112 34
rect 118 29 120 33
rect 150 32 152 46
rect 17 19 19 23
rect 47 19 49 23
rect 55 19 57 23
rect 288 44 290 51
rect 265 37 267 40
rect 824 42 841 44
rect 861 42 874 44
rect 894 42 897 44
rect 824 34 841 36
rect 861 34 874 36
rect 894 34 897 36
rect 288 31 290 34
rect 150 19 152 22
rect 110 15 112 19
rect 118 15 120 19
rect 241 12 243 26
rect 241 -1 243 2
rect 108 -56 110 -52
rect 343 -53 345 -50
rect 15 -72 17 -68
rect 23 -72 25 -68
rect 45 -72 47 -68
rect 53 -72 55 -68
rect 85 -69 87 -65
rect 148 -72 150 -68
rect 15 -105 17 -92
rect 23 -96 25 -92
rect 45 -105 47 -92
rect 53 -105 55 -92
rect 85 -93 87 -89
rect 108 -95 110 -76
rect 920 -55 937 -53
rect 957 -55 970 -53
rect 990 -55 993 -53
rect 920 -63 937 -61
rect 957 -63 970 -61
rect 990 -63 993 -61
rect 231 -78 248 -76
rect 268 -78 281 -76
rect 301 -78 304 -76
rect 231 -86 248 -84
rect 268 -86 281 -84
rect 301 -86 304 -84
rect 343 -87 345 -73
rect 108 -109 110 -104
rect 116 -109 118 -105
rect 148 -106 150 -92
rect 343 -100 345 -97
rect 15 -119 17 -115
rect 45 -119 47 -115
rect 53 -119 55 -115
rect 148 -119 150 -116
rect 108 -123 110 -119
rect 116 -123 118 -119
rect 108 -197 110 -193
rect 15 -213 17 -209
rect 23 -213 25 -209
rect 45 -213 47 -209
rect 53 -213 55 -209
rect 85 -210 87 -206
rect 265 -200 267 -187
rect 288 -200 290 -196
rect 148 -213 150 -209
rect 15 -246 17 -233
rect 23 -237 25 -233
rect 45 -246 47 -233
rect 53 -246 55 -233
rect 85 -234 87 -230
rect 108 -236 110 -217
rect 821 -219 838 -217
rect 858 -219 871 -217
rect 891 -219 894 -217
rect 265 -233 267 -220
rect 288 -224 290 -220
rect 821 -227 838 -225
rect 858 -227 871 -225
rect 891 -227 894 -225
rect 108 -250 110 -245
rect 116 -250 118 -246
rect 148 -247 150 -233
rect 241 -237 243 -234
rect 15 -260 17 -256
rect 45 -260 47 -256
rect 53 -260 55 -256
rect 288 -239 290 -232
rect 265 -246 267 -243
rect 1007 -240 1024 -238
rect 1044 -240 1057 -238
rect 1087 -240 1090 -238
rect 1007 -248 1024 -246
rect 1044 -248 1057 -246
rect 1087 -248 1090 -246
rect 288 -252 290 -249
rect 1007 -256 1024 -254
rect 1044 -256 1057 -254
rect 1087 -256 1090 -254
rect 148 -260 150 -257
rect 108 -264 110 -260
rect 116 -264 118 -260
rect 241 -271 243 -257
rect 241 -284 243 -281
rect 815 -285 832 -283
rect 852 -285 865 -283
rect 895 -285 898 -283
rect 815 -293 832 -291
rect 852 -293 865 -291
rect 895 -293 898 -291
rect 815 -301 832 -299
rect 852 -301 865 -299
rect 895 -301 898 -299
rect 108 -339 110 -335
rect 15 -355 17 -351
rect 23 -355 25 -351
rect 45 -355 47 -351
rect 53 -355 55 -351
rect 85 -352 87 -348
rect 346 -341 348 -338
rect 148 -355 150 -351
rect 15 -388 17 -375
rect 23 -379 25 -375
rect 45 -388 47 -375
rect 53 -388 55 -375
rect 85 -376 87 -372
rect 108 -378 110 -359
rect 231 -361 248 -359
rect 268 -361 281 -359
rect 301 -361 304 -359
rect 231 -369 248 -367
rect 268 -369 281 -367
rect 301 -369 304 -367
rect 346 -375 348 -361
rect 108 -392 110 -387
rect 116 -392 118 -388
rect 148 -389 150 -375
rect 346 -388 348 -385
rect 15 -402 17 -398
rect 45 -402 47 -398
rect 53 -402 55 -398
rect 148 -402 150 -399
rect 108 -406 110 -402
rect 116 -406 118 -402
rect 829 -493 846 -491
rect 866 -493 879 -491
rect 899 -493 902 -491
rect 829 -501 846 -499
rect 866 -501 879 -499
rect 899 -501 902 -499
rect 108 -526 110 -522
rect 15 -542 17 -538
rect 23 -542 25 -538
rect 45 -542 47 -538
rect 53 -542 55 -538
rect 85 -539 87 -535
rect 265 -529 267 -516
rect 288 -529 290 -525
rect 148 -542 150 -538
rect 15 -575 17 -562
rect 23 -566 25 -562
rect 45 -575 47 -562
rect 53 -575 55 -562
rect 85 -563 87 -559
rect 108 -565 110 -546
rect 265 -562 267 -549
rect 288 -553 290 -549
rect 823 -559 840 -557
rect 860 -559 873 -557
rect 903 -559 906 -557
rect 108 -579 110 -574
rect 116 -579 118 -575
rect 148 -576 150 -562
rect 241 -566 243 -563
rect 15 -589 17 -585
rect 45 -589 47 -585
rect 53 -589 55 -585
rect 288 -568 290 -561
rect 823 -567 840 -565
rect 860 -567 873 -565
rect 903 -567 906 -565
rect 265 -575 267 -572
rect 1016 -571 1033 -569
rect 1053 -571 1066 -569
rect 1106 -571 1109 -569
rect 823 -575 840 -573
rect 860 -575 873 -573
rect 903 -575 906 -573
rect 288 -581 290 -578
rect 1016 -579 1033 -577
rect 1053 -579 1066 -577
rect 1106 -579 1109 -577
rect 148 -589 150 -586
rect 108 -593 110 -589
rect 116 -593 118 -589
rect 241 -600 243 -586
rect 1016 -587 1033 -585
rect 1053 -587 1066 -585
rect 1106 -587 1109 -585
rect 1016 -595 1033 -593
rect 1053 -595 1066 -593
rect 1106 -595 1109 -593
rect 241 -613 243 -610
rect 823 -641 840 -639
rect 860 -641 873 -639
rect 913 -641 916 -639
rect 823 -649 840 -647
rect 860 -649 873 -647
rect 913 -649 916 -647
rect 823 -657 840 -655
rect 860 -657 873 -655
rect 913 -657 916 -655
rect 108 -668 110 -664
rect 346 -667 348 -664
rect 823 -665 840 -663
rect 860 -665 873 -663
rect 913 -665 916 -663
rect 15 -684 17 -680
rect 23 -684 25 -680
rect 45 -684 47 -680
rect 53 -684 55 -680
rect 85 -681 87 -677
rect 148 -684 150 -680
rect 15 -717 17 -704
rect 23 -708 25 -704
rect 45 -717 47 -704
rect 53 -717 55 -704
rect 85 -705 87 -701
rect 108 -707 110 -688
rect 231 -690 248 -688
rect 268 -690 281 -688
rect 301 -690 304 -688
rect 231 -698 248 -696
rect 268 -698 281 -696
rect 301 -698 304 -696
rect 346 -701 348 -687
rect 108 -721 110 -716
rect 116 -721 118 -717
rect 148 -718 150 -704
rect 346 -714 348 -711
rect 15 -731 17 -727
rect 45 -731 47 -727
rect 53 -731 55 -727
rect 148 -731 150 -728
rect 108 -735 110 -731
rect 116 -735 118 -731
rect 831 -907 848 -905
rect 868 -907 881 -905
rect 901 -907 904 -905
rect 831 -915 848 -913
rect 868 -915 881 -913
rect 901 -915 904 -913
rect 825 -973 842 -971
rect 862 -973 875 -971
rect 905 -973 908 -971
rect 825 -981 842 -979
rect 862 -981 875 -979
rect 905 -981 908 -979
rect 825 -989 842 -987
rect 862 -989 875 -987
rect 905 -989 908 -987
rect 108 -1016 110 -1012
rect 15 -1032 17 -1028
rect 23 -1032 25 -1028
rect 45 -1032 47 -1028
rect 53 -1032 55 -1028
rect 85 -1029 87 -1025
rect 263 -1018 265 -1005
rect 286 -1018 288 -1014
rect 148 -1032 150 -1028
rect 15 -1065 17 -1052
rect 23 -1056 25 -1052
rect 45 -1065 47 -1052
rect 53 -1065 55 -1052
rect 85 -1053 87 -1049
rect 108 -1055 110 -1036
rect 1041 -1026 1064 -1024
rect 1078 -1026 1091 -1024
rect 1141 -1026 1144 -1024
rect 1041 -1034 1064 -1032
rect 1078 -1034 1091 -1032
rect 1141 -1034 1144 -1032
rect 263 -1051 265 -1038
rect 286 -1042 288 -1038
rect 1041 -1042 1064 -1040
rect 1078 -1042 1091 -1040
rect 1141 -1042 1144 -1040
rect 108 -1069 110 -1064
rect 116 -1069 118 -1065
rect 148 -1066 150 -1052
rect 239 -1055 241 -1052
rect 15 -1079 17 -1075
rect 45 -1079 47 -1075
rect 53 -1079 55 -1075
rect 286 -1057 288 -1050
rect 1041 -1050 1064 -1048
rect 1078 -1050 1091 -1048
rect 1141 -1050 1144 -1048
rect 825 -1055 842 -1053
rect 862 -1055 875 -1053
rect 915 -1055 918 -1053
rect 263 -1064 265 -1061
rect 1041 -1058 1064 -1056
rect 1078 -1058 1091 -1056
rect 1141 -1058 1144 -1056
rect 825 -1063 842 -1061
rect 862 -1063 875 -1061
rect 915 -1063 918 -1061
rect 286 -1070 288 -1067
rect 825 -1071 842 -1069
rect 862 -1071 875 -1069
rect 915 -1071 918 -1069
rect 148 -1079 150 -1076
rect 108 -1083 110 -1079
rect 116 -1083 118 -1079
rect 239 -1089 241 -1075
rect 825 -1079 842 -1077
rect 862 -1079 875 -1077
rect 915 -1079 918 -1077
rect 239 -1102 241 -1099
rect 826 -1142 849 -1140
rect 863 -1142 876 -1140
rect 926 -1142 929 -1140
rect 345 -1152 347 -1149
rect 826 -1150 849 -1148
rect 863 -1150 876 -1148
rect 926 -1150 929 -1148
rect 106 -1157 108 -1153
rect 13 -1173 15 -1169
rect 21 -1173 23 -1169
rect 43 -1173 45 -1169
rect 51 -1173 53 -1169
rect 83 -1170 85 -1166
rect 146 -1173 148 -1169
rect 826 -1158 849 -1156
rect 863 -1158 876 -1156
rect 926 -1158 929 -1156
rect 826 -1166 849 -1164
rect 863 -1166 876 -1164
rect 926 -1166 929 -1164
rect 13 -1206 15 -1193
rect 21 -1197 23 -1193
rect 43 -1206 45 -1193
rect 51 -1206 53 -1193
rect 83 -1194 85 -1190
rect 106 -1196 108 -1177
rect 229 -1179 246 -1177
rect 266 -1179 279 -1177
rect 299 -1179 302 -1177
rect 229 -1187 246 -1185
rect 266 -1187 279 -1185
rect 299 -1187 302 -1185
rect 345 -1186 347 -1172
rect 826 -1174 849 -1172
rect 863 -1174 876 -1172
rect 926 -1174 929 -1172
rect 106 -1210 108 -1205
rect 114 -1210 116 -1206
rect 146 -1207 148 -1193
rect 345 -1199 347 -1196
rect 13 -1220 15 -1216
rect 43 -1220 45 -1216
rect 51 -1220 53 -1216
rect 146 -1220 148 -1217
rect 106 -1224 108 -1220
rect 114 -1224 116 -1220
rect 830 -1402 847 -1400
rect 867 -1402 880 -1400
rect 900 -1402 903 -1400
rect 830 -1410 847 -1408
rect 867 -1410 880 -1408
rect 900 -1410 903 -1408
rect 824 -1468 841 -1466
rect 861 -1468 874 -1466
rect 904 -1468 907 -1466
rect 824 -1476 841 -1474
rect 861 -1476 874 -1474
rect 904 -1476 907 -1474
rect 824 -1484 841 -1482
rect 861 -1484 874 -1482
rect 904 -1484 907 -1482
rect 106 -1506 108 -1502
rect 13 -1522 15 -1518
rect 21 -1522 23 -1518
rect 43 -1522 45 -1518
rect 51 -1522 53 -1518
rect 83 -1519 85 -1515
rect 262 -1508 264 -1495
rect 285 -1508 287 -1504
rect 146 -1522 148 -1518
rect 13 -1555 15 -1542
rect 21 -1546 23 -1542
rect 43 -1555 45 -1542
rect 51 -1555 53 -1542
rect 83 -1543 85 -1539
rect 106 -1545 108 -1526
rect 262 -1541 264 -1528
rect 285 -1532 287 -1528
rect 1048 -1534 1065 -1532
rect 1085 -1534 1098 -1532
rect 1158 -1534 1161 -1532
rect 106 -1559 108 -1554
rect 114 -1559 116 -1555
rect 146 -1556 148 -1542
rect 238 -1545 240 -1542
rect 13 -1569 15 -1565
rect 43 -1569 45 -1565
rect 51 -1569 53 -1565
rect 285 -1547 287 -1540
rect 1048 -1542 1065 -1540
rect 1085 -1542 1098 -1540
rect 1158 -1542 1161 -1540
rect 262 -1554 264 -1551
rect 824 -1550 841 -1548
rect 861 -1550 874 -1548
rect 914 -1550 917 -1548
rect 1048 -1550 1065 -1548
rect 1085 -1550 1098 -1548
rect 1158 -1550 1161 -1548
rect 285 -1560 287 -1557
rect 824 -1558 841 -1556
rect 861 -1558 874 -1556
rect 914 -1558 917 -1556
rect 1048 -1558 1065 -1556
rect 1085 -1558 1098 -1556
rect 1158 -1558 1161 -1556
rect 146 -1569 148 -1566
rect 106 -1573 108 -1569
rect 114 -1573 116 -1569
rect 238 -1579 240 -1565
rect 824 -1566 841 -1564
rect 861 -1566 874 -1564
rect 914 -1566 917 -1564
rect 1048 -1566 1065 -1564
rect 1085 -1566 1098 -1564
rect 1158 -1566 1161 -1564
rect 824 -1574 841 -1572
rect 861 -1574 874 -1572
rect 914 -1574 917 -1572
rect 1048 -1574 1065 -1572
rect 1085 -1574 1098 -1572
rect 1158 -1574 1161 -1572
rect 238 -1592 240 -1589
rect 345 -1638 347 -1635
rect 825 -1637 848 -1635
rect 862 -1637 875 -1635
rect 925 -1637 928 -1635
rect 106 -1647 108 -1643
rect 13 -1663 15 -1659
rect 21 -1663 23 -1659
rect 43 -1663 45 -1659
rect 51 -1663 53 -1659
rect 83 -1660 85 -1656
rect 825 -1645 848 -1643
rect 862 -1645 875 -1643
rect 925 -1645 928 -1643
rect 825 -1653 848 -1651
rect 862 -1653 875 -1651
rect 925 -1653 928 -1651
rect 146 -1663 148 -1659
rect 13 -1696 15 -1683
rect 21 -1687 23 -1683
rect 43 -1696 45 -1683
rect 51 -1696 53 -1683
rect 83 -1684 85 -1680
rect 106 -1686 108 -1667
rect 228 -1669 245 -1667
rect 265 -1669 278 -1667
rect 298 -1669 301 -1667
rect 345 -1672 347 -1658
rect 825 -1661 848 -1659
rect 862 -1661 875 -1659
rect 925 -1661 928 -1659
rect 825 -1669 848 -1667
rect 862 -1669 875 -1667
rect 925 -1669 928 -1667
rect 228 -1677 245 -1675
rect 265 -1677 278 -1675
rect 298 -1677 301 -1675
rect 106 -1700 108 -1695
rect 114 -1700 116 -1696
rect 146 -1697 148 -1683
rect 345 -1685 347 -1682
rect 13 -1710 15 -1706
rect 43 -1710 45 -1706
rect 51 -1710 53 -1706
rect 146 -1710 148 -1707
rect 106 -1714 108 -1710
rect 114 -1714 116 -1710
rect 821 -1741 838 -1739
rect 858 -1741 871 -1739
rect 931 -1741 934 -1739
rect 821 -1749 838 -1747
rect 858 -1749 871 -1747
rect 931 -1749 934 -1747
rect 821 -1757 838 -1755
rect 858 -1757 871 -1755
rect 931 -1757 934 -1755
rect 821 -1765 838 -1763
rect 858 -1765 871 -1763
rect 931 -1765 934 -1763
rect 821 -1773 838 -1771
rect 858 -1773 871 -1771
rect 931 -1773 934 -1771
rect 821 -1781 838 -1779
rect 858 -1781 871 -1779
rect 931 -1781 934 -1779
rect 106 -1976 108 -1972
rect 13 -1992 15 -1988
rect 21 -1992 23 -1988
rect 43 -1992 45 -1988
rect 51 -1992 53 -1988
rect 83 -1989 85 -1985
rect 146 -1992 148 -1988
rect 13 -2025 15 -2012
rect 21 -2016 23 -2012
rect 43 -2025 45 -2012
rect 51 -2025 53 -2012
rect 83 -2013 85 -2009
rect 106 -2015 108 -1996
rect 106 -2029 108 -2024
rect 114 -2029 116 -2025
rect 146 -2026 148 -2012
rect 13 -2039 15 -2035
rect 43 -2039 45 -2035
rect 51 -2039 53 -2035
rect 146 -2039 148 -2036
rect 106 -2043 108 -2039
rect 114 -2043 116 -2039
<< polycontact >>
rect 265 96 269 100
rect 285 87 290 92
rect 17 70 21 74
rect 54 70 58 74
rect 87 73 91 77
rect 106 55 110 59
rect 106 43 110 47
rect 106 32 110 36
rect 146 35 150 39
rect 820 42 824 46
rect 820 34 824 38
rect 288 27 292 31
rect 237 15 241 19
rect 15 -68 19 -64
rect 52 -68 56 -64
rect 85 -65 89 -61
rect 104 -83 108 -79
rect 104 -95 108 -91
rect 227 -78 231 -74
rect 916 -55 920 -51
rect 916 -63 920 -59
rect 227 -86 231 -82
rect 339 -84 343 -80
rect 104 -106 108 -102
rect 144 -103 148 -99
rect 265 -187 269 -183
rect 15 -209 19 -205
rect 52 -209 56 -205
rect 85 -206 89 -202
rect 285 -196 290 -191
rect 104 -224 108 -220
rect 104 -236 108 -232
rect 817 -219 821 -215
rect 817 -227 821 -223
rect 104 -247 108 -243
rect 144 -244 148 -240
rect 1003 -240 1007 -236
rect 1003 -248 1007 -244
rect 288 -256 292 -252
rect 1003 -256 1007 -252
rect 237 -268 241 -264
rect 811 -285 815 -281
rect 811 -293 815 -289
rect 811 -301 815 -297
rect 15 -351 19 -347
rect 52 -351 56 -347
rect 85 -348 89 -344
rect 104 -366 108 -362
rect 104 -378 108 -374
rect 227 -361 231 -357
rect 227 -369 231 -365
rect 342 -372 346 -368
rect 104 -389 108 -385
rect 144 -386 148 -382
rect 825 -493 829 -489
rect 825 -501 829 -497
rect 265 -516 269 -512
rect 15 -538 19 -534
rect 52 -538 56 -534
rect 85 -535 89 -531
rect 285 -525 290 -520
rect 104 -553 108 -549
rect 104 -565 108 -561
rect 819 -559 823 -555
rect 104 -576 108 -572
rect 144 -573 148 -569
rect 819 -567 823 -563
rect 819 -575 823 -571
rect 1012 -571 1016 -567
rect 1012 -579 1016 -575
rect 288 -585 292 -581
rect 237 -597 241 -593
rect 1012 -587 1016 -583
rect 1012 -595 1016 -591
rect 819 -641 823 -637
rect 819 -649 823 -645
rect 819 -657 823 -653
rect 819 -665 823 -661
rect 15 -680 19 -676
rect 52 -680 56 -676
rect 85 -677 89 -673
rect 104 -695 108 -691
rect 104 -707 108 -703
rect 227 -690 231 -686
rect 227 -698 231 -694
rect 342 -698 346 -694
rect 104 -718 108 -714
rect 144 -715 148 -711
rect 827 -907 831 -903
rect 827 -915 831 -911
rect 821 -973 825 -969
rect 821 -981 825 -977
rect 821 -989 825 -985
rect 263 -1005 267 -1001
rect 15 -1028 19 -1024
rect 52 -1028 56 -1024
rect 85 -1025 89 -1021
rect 283 -1014 288 -1009
rect 104 -1043 108 -1039
rect 104 -1055 108 -1051
rect 1037 -1027 1041 -1023
rect 1037 -1035 1041 -1031
rect 1037 -1043 1041 -1039
rect 104 -1066 108 -1062
rect 144 -1063 148 -1059
rect 821 -1055 825 -1051
rect 1037 -1051 1041 -1047
rect 821 -1063 825 -1059
rect 1037 -1059 1041 -1055
rect 286 -1074 290 -1070
rect 821 -1071 825 -1067
rect 235 -1086 239 -1082
rect 821 -1079 825 -1075
rect 822 -1143 826 -1139
rect 822 -1151 826 -1147
rect 13 -1169 17 -1165
rect 50 -1169 54 -1165
rect 83 -1166 87 -1162
rect 822 -1159 826 -1155
rect 822 -1167 826 -1163
rect 102 -1184 106 -1180
rect 102 -1196 106 -1192
rect 225 -1179 229 -1175
rect 225 -1187 229 -1183
rect 341 -1183 345 -1179
rect 822 -1177 826 -1172
rect 102 -1207 106 -1203
rect 142 -1204 146 -1200
rect 826 -1402 830 -1398
rect 826 -1410 830 -1406
rect 820 -1468 824 -1464
rect 820 -1476 824 -1472
rect 820 -1484 824 -1480
rect 262 -1495 266 -1491
rect 13 -1518 17 -1514
rect 50 -1518 54 -1514
rect 83 -1515 87 -1511
rect 282 -1504 287 -1499
rect 102 -1533 106 -1529
rect 102 -1545 106 -1541
rect 1044 -1534 1048 -1530
rect 102 -1556 106 -1552
rect 142 -1553 146 -1549
rect 1044 -1542 1048 -1538
rect 820 -1550 824 -1546
rect 1044 -1550 1048 -1546
rect 820 -1558 824 -1554
rect 1044 -1558 1048 -1554
rect 285 -1564 289 -1560
rect 234 -1576 238 -1572
rect 820 -1566 824 -1562
rect 1044 -1566 1048 -1562
rect 820 -1574 824 -1570
rect 1044 -1574 1048 -1570
rect 821 -1638 825 -1634
rect 13 -1659 17 -1655
rect 50 -1659 54 -1655
rect 83 -1656 87 -1652
rect 821 -1646 825 -1642
rect 821 -1654 825 -1650
rect 102 -1674 106 -1670
rect 102 -1686 106 -1682
rect 224 -1669 228 -1665
rect 341 -1669 345 -1665
rect 224 -1677 228 -1673
rect 821 -1662 825 -1658
rect 821 -1671 825 -1667
rect 102 -1697 106 -1693
rect 142 -1694 146 -1690
rect 817 -1741 821 -1737
rect 817 -1749 821 -1745
rect 817 -1757 821 -1753
rect 817 -1765 821 -1761
rect 817 -1774 821 -1770
rect 817 -1783 821 -1779
rect 13 -1988 17 -1984
rect 50 -1988 54 -1984
rect 83 -1985 87 -1981
rect 102 -2003 106 -1999
rect 102 -2015 106 -2011
rect 102 -2026 106 -2022
rect 142 -2023 146 -2019
<< metal1 >>
rect -17 128 523 131
rect -17 0 -14 128
rect 207 108 269 112
rect 9 90 155 94
rect 159 90 162 94
rect 9 62 12 90
rect 17 74 21 77
rect 39 62 42 90
rect 50 82 61 87
rect 54 74 59 82
rect 58 70 59 74
rect 79 62 82 90
rect 105 82 109 90
rect 87 77 91 80
rect 94 66 100 69
rect 97 59 100 66
rect 97 55 106 59
rect 28 43 32 46
rect 58 42 62 46
rect 101 43 106 47
rect 101 42 105 43
rect 58 38 105 42
rect 28 33 32 38
rect 58 33 62 38
rect 101 36 105 38
rect 121 39 125 62
rect 145 66 149 90
rect 153 39 157 46
rect 207 39 211 108
rect 265 101 269 108
rect 265 100 308 101
rect 269 96 308 100
rect 260 87 285 92
rect 225 83 264 87
rect 225 70 229 83
rect 226 63 229 70
rect 101 32 106 36
rect 121 35 146 39
rect 153 35 211 39
rect 121 29 125 35
rect 153 32 157 35
rect 12 5 16 23
rect 42 5 47 23
rect 105 5 109 19
rect 145 5 149 22
rect 225 19 229 63
rect 237 54 241 59
rect 268 57 272 63
rect 283 57 287 63
rect 268 53 287 57
rect 268 50 272 53
rect 236 46 240 50
rect 244 19 248 26
rect 275 46 279 53
rect 283 44 287 53
rect 260 19 264 40
rect 291 57 295 63
rect 303 57 308 96
rect 291 53 308 57
rect 291 44 295 53
rect 391 37 395 104
rect 399 48 403 104
rect 288 19 292 27
rect 225 15 237 19
rect 244 15 292 19
rect 244 12 248 15
rect -4 0 0 5
rect 4 0 224 5
rect -19 -6 2 0
rect 219 -1 224 0
rect 236 -1 240 2
rect 219 -2 240 -1
rect 219 -6 236 -2
rect -4 -133 2 -6
rect 7 -48 153 -44
rect 157 -48 160 -44
rect 7 -76 10 -48
rect 15 -64 19 -61
rect 37 -76 40 -48
rect 48 -56 59 -51
rect 52 -64 57 -56
rect 56 -68 57 -64
rect 77 -76 80 -48
rect 103 -56 107 -48
rect 92 -72 98 -69
rect 95 -79 98 -72
rect 95 -83 104 -79
rect 26 -95 30 -92
rect 56 -96 60 -92
rect 99 -95 104 -91
rect 99 -96 103 -95
rect 56 -100 103 -96
rect 26 -105 30 -100
rect 56 -105 60 -100
rect 99 -102 103 -100
rect 119 -99 123 -76
rect 143 -72 147 -48
rect 338 -53 342 -49
rect 274 -66 325 -62
rect 274 -71 278 -66
rect 151 -99 155 -92
rect 239 -75 248 -71
rect 274 -75 281 -71
rect 168 -86 227 -82
rect 168 -99 172 -86
rect 239 -87 243 -75
rect 274 -79 278 -75
rect 268 -83 278 -79
rect 321 -80 325 -66
rect 346 -80 350 -73
rect 321 -84 339 -80
rect 346 -84 356 -80
rect 243 -91 248 -87
rect 301 -91 305 -87
rect 346 -87 350 -84
rect 99 -106 104 -102
rect 119 -103 144 -99
rect 151 -103 172 -99
rect 119 -109 123 -103
rect 151 -106 155 -103
rect 10 -133 14 -115
rect 40 -133 45 -115
rect 103 -133 107 -119
rect 143 -133 147 -116
rect 305 -133 309 -91
rect 338 -101 342 -97
rect 338 -133 342 -105
rect -4 -138 -2 -133
rect 2 -138 342 -133
rect -4 -274 2 -138
rect 209 -177 269 -173
rect 7 -189 153 -185
rect 157 -189 160 -185
rect 7 -217 10 -189
rect 15 -205 19 -202
rect 37 -217 40 -189
rect 48 -197 59 -192
rect 52 -205 57 -197
rect 56 -209 57 -205
rect 77 -217 80 -189
rect 103 -197 107 -189
rect 92 -213 98 -210
rect 95 -220 98 -213
rect 95 -224 104 -220
rect 26 -236 30 -233
rect 56 -237 60 -233
rect 99 -236 104 -232
rect 99 -237 103 -236
rect 56 -241 103 -237
rect 26 -246 30 -241
rect 56 -246 60 -241
rect 99 -243 103 -241
rect 119 -240 123 -217
rect 143 -213 147 -189
rect 151 -240 155 -233
rect 209 -239 213 -177
rect 265 -182 269 -177
rect 265 -183 308 -182
rect 269 -187 308 -183
rect 260 -196 285 -191
rect 225 -200 264 -196
rect 99 -247 104 -243
rect 119 -244 144 -240
rect 151 -244 209 -240
rect 119 -250 123 -244
rect 151 -247 155 -244
rect 10 -274 14 -256
rect 40 -274 45 -256
rect 103 -274 107 -260
rect 143 -274 147 -257
rect 225 -264 229 -200
rect 237 -229 241 -224
rect 268 -226 272 -220
rect 283 -226 287 -220
rect 268 -230 287 -226
rect 268 -233 272 -230
rect 236 -237 240 -233
rect 244 -264 248 -257
rect 275 -237 279 -230
rect 283 -239 287 -230
rect 260 -264 264 -243
rect 291 -226 295 -220
rect 303 -226 308 -187
rect 291 -230 308 -226
rect 291 -239 295 -230
rect 288 -264 292 -256
rect 225 -268 237 -264
rect 244 -268 292 -264
rect 244 -271 248 -268
rect -4 -279 -2 -274
rect 2 -279 216 -274
rect -4 -416 2 -279
rect 211 -284 216 -279
rect 236 -284 240 -281
rect 211 -285 240 -284
rect 211 -289 236 -285
rect 391 -297 395 32
rect 399 11 403 43
rect 399 -288 403 6
rect 407 -80 411 104
rect 407 -224 411 -85
rect 415 -59 419 104
rect 415 -89 419 -64
rect 7 -331 153 -327
rect 157 -331 160 -327
rect 7 -359 10 -331
rect 15 -347 19 -344
rect 37 -359 40 -331
rect 48 -339 59 -334
rect 52 -347 57 -339
rect 56 -351 57 -347
rect 77 -359 80 -331
rect 103 -339 107 -331
rect 92 -355 98 -352
rect 95 -362 98 -355
rect 95 -366 104 -362
rect 26 -378 30 -375
rect 56 -379 60 -375
rect 99 -378 104 -374
rect 99 -379 103 -378
rect 56 -383 103 -379
rect 26 -388 30 -383
rect 56 -388 60 -383
rect 99 -385 103 -383
rect 119 -382 123 -359
rect 143 -355 147 -331
rect 341 -341 345 -337
rect 274 -345 326 -341
rect 274 -354 278 -345
rect 225 -361 227 -357
rect 239 -358 248 -354
rect 274 -358 281 -354
rect 151 -382 155 -375
rect 180 -368 227 -365
rect 175 -369 227 -368
rect 175 -382 179 -369
rect 239 -370 243 -358
rect 274 -362 278 -358
rect 268 -366 278 -362
rect 322 -368 326 -345
rect 349 -368 353 -361
rect 243 -374 248 -370
rect 301 -374 305 -370
rect 322 -372 342 -368
rect 349 -372 363 -368
rect 99 -389 104 -385
rect 119 -386 144 -382
rect 151 -386 179 -382
rect 119 -392 123 -386
rect 151 -389 155 -386
rect 10 -416 14 -398
rect 40 -416 45 -398
rect 103 -416 107 -402
rect 143 -416 147 -399
rect 305 -416 310 -374
rect 349 -375 353 -372
rect 341 -389 345 -385
rect 340 -416 345 -393
rect -4 -421 -2 -416
rect 2 -421 345 -416
rect -4 -603 2 -421
rect 207 -505 269 -501
rect 7 -518 153 -514
rect 157 -518 160 -514
rect 7 -546 10 -518
rect 15 -534 19 -531
rect 37 -546 40 -518
rect 48 -526 59 -521
rect 52 -534 57 -526
rect 56 -538 57 -534
rect 77 -546 80 -518
rect 103 -526 107 -518
rect 92 -542 98 -539
rect 95 -549 98 -542
rect 95 -553 104 -549
rect 26 -565 30 -562
rect 56 -566 60 -562
rect 99 -565 104 -561
rect 99 -566 103 -565
rect 56 -570 103 -566
rect 26 -575 30 -570
rect 56 -575 60 -570
rect 99 -572 103 -570
rect 119 -569 123 -546
rect 143 -542 147 -518
rect 151 -569 155 -562
rect 207 -568 211 -505
rect 265 -511 269 -505
rect 265 -512 308 -511
rect 269 -516 308 -512
rect 260 -525 285 -520
rect 225 -529 264 -525
rect 99 -576 104 -572
rect 119 -573 144 -569
rect 151 -573 207 -569
rect 119 -579 123 -573
rect 151 -576 155 -573
rect 10 -603 14 -585
rect 40 -603 45 -585
rect 103 -603 107 -589
rect 143 -603 147 -586
rect 225 -593 229 -529
rect 237 -558 241 -553
rect 268 -555 272 -549
rect 283 -555 287 -549
rect 268 -559 287 -555
rect 268 -562 272 -559
rect 236 -566 240 -562
rect 244 -593 248 -586
rect 275 -566 279 -559
rect 283 -568 287 -559
rect 260 -593 264 -572
rect 291 -555 295 -549
rect 303 -555 308 -516
rect 291 -559 308 -555
rect 291 -568 295 -559
rect 288 -593 292 -585
rect 225 -597 237 -593
rect 244 -597 292 -593
rect 244 -600 248 -597
rect -4 -608 -2 -603
rect 2 -608 215 -603
rect -4 -745 2 -608
rect 210 -613 215 -608
rect 236 -613 240 -610
rect 210 -614 240 -613
rect 210 -618 236 -614
rect 7 -660 153 -656
rect 157 -660 160 -656
rect 7 -688 10 -660
rect 15 -676 19 -673
rect 37 -688 40 -660
rect 48 -668 59 -663
rect 52 -676 57 -668
rect 56 -680 57 -676
rect 77 -688 80 -660
rect 103 -668 107 -660
rect 92 -684 98 -681
rect 95 -691 98 -684
rect 95 -695 104 -691
rect 26 -707 30 -704
rect 56 -708 60 -704
rect 99 -707 104 -703
rect 99 -708 103 -707
rect 56 -712 103 -708
rect 26 -717 30 -712
rect 56 -717 60 -712
rect 99 -714 103 -712
rect 119 -711 123 -688
rect 143 -684 147 -660
rect 341 -667 345 -663
rect 391 -663 395 -302
rect 399 -654 403 -293
rect 407 -572 411 -229
rect 274 -674 325 -670
rect 274 -683 278 -674
rect 226 -690 227 -686
rect 239 -687 248 -683
rect 274 -687 281 -683
rect 151 -711 155 -704
rect 208 -698 227 -694
rect 99 -718 104 -714
rect 119 -715 144 -711
rect 151 -715 170 -711
rect 208 -711 212 -698
rect 239 -699 243 -687
rect 274 -691 278 -687
rect 268 -695 278 -691
rect 321 -694 325 -674
rect 349 -694 353 -687
rect 321 -698 342 -694
rect 349 -698 363 -694
rect 243 -703 248 -699
rect 301 -703 305 -699
rect 349 -701 353 -698
rect 177 -715 212 -711
rect 119 -721 123 -715
rect 151 -718 155 -715
rect 10 -745 14 -727
rect 40 -745 45 -727
rect 103 -745 107 -731
rect 143 -745 147 -728
rect 305 -745 310 -703
rect 341 -715 345 -711
rect 340 -745 345 -719
rect -4 -750 -2 -745
rect 2 -750 345 -745
rect -4 -1093 2 -750
rect 208 -995 267 -991
rect 7 -1008 153 -1004
rect 157 -1008 160 -1004
rect 7 -1036 10 -1008
rect 15 -1024 19 -1021
rect 37 -1036 40 -1008
rect 48 -1016 59 -1011
rect 52 -1024 57 -1016
rect 56 -1028 57 -1024
rect 77 -1036 80 -1008
rect 103 -1016 107 -1008
rect 92 -1032 98 -1029
rect 95 -1039 98 -1032
rect 95 -1043 104 -1039
rect 26 -1055 30 -1052
rect 56 -1056 60 -1052
rect 99 -1055 104 -1051
rect 99 -1056 103 -1055
rect 56 -1060 103 -1056
rect 26 -1065 30 -1060
rect 56 -1065 60 -1060
rect 99 -1062 103 -1060
rect 119 -1059 123 -1036
rect 143 -1032 147 -1008
rect 151 -1059 155 -1052
rect 208 -1059 212 -995
rect 263 -1000 267 -995
rect 263 -1001 306 -1000
rect 267 -1005 306 -1001
rect 258 -1014 283 -1009
rect 223 -1018 262 -1014
rect 223 -1042 227 -1018
rect 223 -1047 229 -1042
rect 237 -1047 241 -1042
rect 266 -1044 270 -1038
rect 281 -1044 285 -1038
rect 99 -1066 104 -1062
rect 119 -1063 144 -1059
rect 151 -1063 208 -1059
rect 119 -1069 123 -1063
rect 151 -1066 155 -1063
rect 10 -1093 14 -1075
rect 40 -1093 45 -1075
rect 103 -1093 107 -1079
rect 143 -1093 147 -1076
rect 223 -1082 227 -1047
rect 266 -1048 285 -1044
rect 266 -1051 270 -1048
rect 234 -1055 238 -1051
rect 242 -1082 246 -1075
rect 273 -1055 277 -1048
rect 281 -1057 285 -1048
rect 258 -1082 262 -1061
rect 289 -1044 293 -1038
rect 301 -1044 306 -1005
rect 289 -1048 306 -1044
rect 289 -1057 293 -1048
rect 286 -1082 290 -1074
rect 223 -1086 235 -1082
rect 242 -1086 290 -1082
rect 242 -1089 246 -1086
rect -4 -1098 -2 -1093
rect 2 -1098 209 -1093
rect -4 -1234 2 -1098
rect 204 -1102 209 -1098
rect 234 -1102 238 -1099
rect 204 -1103 238 -1102
rect 204 -1107 234 -1103
rect 5 -1149 151 -1145
rect 155 -1149 158 -1145
rect 5 -1177 8 -1149
rect 13 -1165 17 -1162
rect 35 -1177 38 -1149
rect 46 -1157 57 -1152
rect 50 -1165 55 -1157
rect 54 -1169 55 -1165
rect 75 -1177 78 -1149
rect 101 -1157 105 -1149
rect 90 -1173 96 -1170
rect 93 -1180 96 -1173
rect 93 -1184 102 -1180
rect 24 -1196 28 -1193
rect 54 -1197 58 -1193
rect 97 -1196 102 -1192
rect 97 -1197 101 -1196
rect 54 -1201 101 -1197
rect 24 -1206 28 -1201
rect 54 -1206 58 -1201
rect 97 -1203 101 -1201
rect 117 -1200 121 -1177
rect 141 -1173 145 -1149
rect 340 -1152 344 -1148
rect 391 -1152 395 -668
rect 272 -1163 317 -1159
rect 272 -1172 276 -1163
rect 218 -1179 225 -1175
rect 237 -1176 246 -1172
rect 272 -1176 279 -1172
rect 149 -1200 153 -1193
rect 178 -1187 225 -1183
rect 173 -1200 177 -1187
rect 237 -1188 241 -1176
rect 272 -1180 276 -1176
rect 313 -1179 317 -1163
rect 348 -1179 352 -1172
rect 266 -1184 276 -1180
rect 313 -1183 341 -1179
rect 348 -1183 362 -1179
rect 348 -1186 352 -1183
rect 241 -1192 246 -1188
rect 299 -1192 303 -1188
rect 97 -1207 102 -1203
rect 117 -1204 142 -1200
rect 149 -1204 177 -1200
rect 117 -1210 121 -1204
rect 149 -1207 153 -1204
rect 8 -1234 12 -1216
rect 38 -1234 43 -1216
rect 101 -1234 105 -1220
rect 141 -1234 145 -1217
rect 302 -1234 307 -1192
rect 340 -1200 344 -1196
rect 339 -1234 344 -1204
rect 0 -1239 344 -1234
rect -4 -1378 2 -1239
rect -9 -1382 2 -1378
rect -4 -1583 2 -1382
rect 196 -1481 266 -1477
rect 5 -1498 151 -1494
rect 155 -1498 158 -1494
rect 5 -1526 8 -1498
rect 13 -1514 17 -1511
rect 35 -1526 38 -1498
rect 46 -1506 57 -1501
rect 50 -1514 55 -1506
rect 54 -1518 55 -1514
rect 75 -1526 78 -1498
rect 101 -1506 105 -1498
rect 83 -1511 88 -1506
rect 90 -1522 96 -1519
rect 93 -1529 96 -1522
rect 93 -1533 102 -1529
rect 24 -1545 28 -1542
rect 54 -1546 58 -1542
rect 97 -1545 102 -1541
rect 97 -1546 101 -1545
rect 54 -1550 101 -1546
rect 24 -1555 28 -1550
rect 54 -1555 58 -1550
rect 97 -1552 101 -1550
rect 117 -1549 121 -1526
rect 141 -1522 145 -1498
rect 149 -1549 153 -1542
rect 196 -1549 200 -1481
rect 262 -1490 266 -1481
rect 262 -1491 305 -1490
rect 266 -1495 305 -1491
rect 257 -1504 282 -1499
rect 222 -1508 261 -1504
rect 222 -1516 226 -1508
rect 223 -1522 226 -1516
rect 222 -1532 226 -1522
rect 222 -1537 229 -1532
rect 237 -1537 241 -1532
rect 265 -1534 269 -1528
rect 280 -1534 284 -1528
rect 97 -1556 102 -1552
rect 117 -1553 142 -1549
rect 149 -1553 196 -1549
rect 117 -1559 121 -1553
rect 149 -1556 153 -1553
rect 8 -1583 12 -1565
rect 38 -1583 43 -1565
rect 101 -1583 105 -1569
rect 141 -1583 145 -1566
rect 222 -1572 226 -1537
rect 265 -1538 284 -1534
rect 265 -1541 269 -1538
rect 233 -1545 237 -1541
rect 241 -1572 245 -1565
rect 272 -1545 276 -1538
rect 280 -1547 284 -1538
rect 257 -1572 261 -1551
rect 288 -1534 292 -1528
rect 300 -1534 305 -1495
rect 288 -1538 305 -1534
rect 288 -1547 292 -1538
rect 285 -1572 289 -1564
rect 222 -1576 234 -1572
rect 241 -1576 289 -1572
rect 241 -1579 245 -1576
rect 0 -1588 205 -1583
rect -4 -1724 2 -1588
rect 200 -1592 205 -1588
rect 233 -1592 237 -1589
rect 200 -1593 237 -1592
rect 200 -1597 233 -1593
rect 5 -1639 151 -1635
rect 155 -1639 158 -1635
rect 340 -1638 344 -1634
rect 5 -1667 8 -1639
rect 13 -1655 17 -1652
rect 35 -1667 38 -1639
rect 46 -1647 57 -1642
rect 50 -1655 55 -1647
rect 54 -1659 55 -1655
rect 75 -1667 78 -1639
rect 101 -1647 105 -1639
rect 90 -1663 96 -1660
rect 93 -1670 96 -1663
rect 93 -1674 102 -1670
rect 24 -1686 28 -1683
rect 54 -1687 58 -1683
rect 97 -1686 102 -1682
rect 97 -1687 101 -1686
rect 54 -1691 101 -1687
rect 24 -1696 28 -1691
rect 54 -1696 58 -1691
rect 97 -1693 101 -1691
rect 117 -1690 121 -1667
rect 141 -1663 145 -1639
rect 271 -1650 326 -1646
rect 271 -1662 275 -1650
rect 222 -1669 224 -1665
rect 236 -1666 245 -1662
rect 271 -1666 278 -1662
rect 322 -1665 326 -1650
rect 348 -1665 352 -1658
rect 149 -1690 153 -1683
rect 181 -1677 224 -1673
rect 176 -1690 180 -1677
rect 236 -1678 240 -1666
rect 271 -1670 275 -1666
rect 322 -1669 341 -1665
rect 348 -1669 362 -1665
rect 265 -1674 275 -1670
rect 348 -1672 352 -1669
rect 240 -1682 245 -1678
rect 298 -1682 302 -1678
rect 97 -1697 102 -1693
rect 117 -1694 142 -1690
rect 149 -1694 180 -1690
rect 117 -1700 121 -1694
rect 149 -1697 153 -1694
rect 8 -1724 12 -1706
rect 38 -1724 43 -1706
rect 101 -1724 105 -1710
rect 141 -1724 145 -1707
rect 302 -1724 307 -1682
rect 340 -1686 344 -1682
rect 339 -1724 344 -1690
rect 0 -1729 344 -1724
rect -4 -2053 2 -1729
rect 391 -1786 395 -1158
rect 399 -1165 403 -659
rect 407 -1077 411 -577
rect 399 -1770 403 -1170
rect 407 -1658 411 -1082
rect 5 -1968 151 -1964
rect 155 -1968 158 -1964
rect 5 -1996 8 -1968
rect 13 -1984 17 -1981
rect 35 -1996 38 -1968
rect 46 -1976 57 -1971
rect 50 -1984 55 -1976
rect 54 -1988 55 -1984
rect 75 -1996 78 -1968
rect 101 -1976 105 -1968
rect 90 -1992 96 -1989
rect 93 -1999 96 -1992
rect 93 -2003 102 -1999
rect 24 -2015 28 -2012
rect 54 -2016 58 -2012
rect 97 -2015 102 -2011
rect 97 -2016 101 -2015
rect 54 -2020 101 -2016
rect 24 -2025 28 -2020
rect 54 -2025 58 -2020
rect 97 -2022 101 -2020
rect 117 -2019 121 -1996
rect 141 -1992 145 -1968
rect 149 -2019 153 -2012
rect 391 -2019 395 -1791
rect 97 -2026 102 -2022
rect 117 -2023 142 -2019
rect 149 -2023 160 -2019
rect 117 -2029 121 -2023
rect 149 -2026 153 -2023
rect 8 -2053 12 -2035
rect 38 -2053 43 -2035
rect 101 -2053 105 -2039
rect 141 -2053 145 -2036
rect 391 -2042 395 -2024
rect 399 -2042 403 -1775
rect 407 -2042 411 -1664
rect 415 -2042 419 -94
rect 423 -213 427 104
rect 423 -271 427 -218
rect 423 -280 427 -276
rect 423 -563 427 -285
rect 431 -368 435 104
rect 431 -499 435 -373
rect 439 -257 443 104
rect 439 -379 443 -263
rect 423 -645 427 -568
rect 423 -1067 427 -650
rect 431 -985 435 -504
rect 423 -1156 427 -1073
rect 423 -1660 427 -1161
rect 431 -1568 435 -991
rect 423 -1769 427 -1665
rect 423 -2042 427 -1774
rect 431 -2042 435 -1573
rect 439 -2042 443 -384
rect 447 -489 451 104
rect 447 -554 451 -494
rect 447 -600 451 -559
rect 447 -636 451 -605
rect 447 -977 451 -641
rect 455 -694 459 104
rect 455 -911 459 -699
rect 463 -604 467 104
rect 463 -704 467 -609
rect 447 -1045 451 -982
rect 447 -1147 451 -1050
rect 447 -1563 451 -1152
rect 455 -1481 459 -916
rect 447 -1651 451 -1568
rect 447 -1760 451 -1656
rect 447 -2042 451 -1765
rect 455 -2042 459 -1486
rect 463 -2042 467 -709
rect 471 -902 475 104
rect 471 -968 475 -907
rect 471 -1032 475 -973
rect 471 -1056 475 -1038
rect 471 -1138 475 -1061
rect 471 -1472 475 -1143
rect 479 -1179 483 104
rect 479 -1407 483 -1184
rect 487 -1020 491 104
rect 487 -1242 491 -1026
rect 471 -1554 475 -1477
rect 471 -1642 475 -1559
rect 471 -1751 475 -1647
rect 471 -2042 475 -1756
rect 479 -2042 483 -1412
rect 487 -2042 491 -1247
rect 495 -1398 499 104
rect 495 -1463 499 -1403
rect 495 -1545 499 -1468
rect 495 -1580 499 -1550
rect 495 -1633 499 -1585
rect 495 -1742 499 -1638
rect 503 -1674 507 104
rect 495 -2042 499 -1747
rect 503 -2042 507 -1679
rect 511 -1733 515 104
rect 511 -2042 515 -1738
rect 519 -2042 523 128
rect 867 59 909 63
rect 867 49 871 59
rect 819 42 820 46
rect 832 45 841 49
rect 867 45 874 49
rect 819 34 820 38
rect 832 33 836 45
rect 867 41 871 45
rect 861 37 871 41
rect 836 29 841 33
rect 894 29 898 33
rect 905 -51 909 59
rect 963 -48 967 -39
rect 905 -55 916 -51
rect 928 -52 937 -48
rect 963 -52 970 -48
rect 914 -63 916 -59
rect 928 -64 932 -52
rect 963 -56 967 -52
rect 957 -60 967 -56
rect 932 -68 937 -64
rect 990 -68 993 -64
rect 864 -207 995 -203
rect 864 -212 868 -207
rect 815 -219 817 -215
rect 829 -216 838 -212
rect 864 -216 871 -212
rect 815 -227 817 -223
rect 829 -228 833 -216
rect 864 -220 868 -216
rect 858 -224 868 -220
rect 833 -232 838 -228
rect 891 -232 894 -228
rect 991 -236 995 -207
rect 1050 -233 1054 -224
rect 991 -240 1003 -236
rect 1044 -237 1057 -233
rect 987 -248 1003 -244
rect 1015 -245 1024 -241
rect 991 -256 1003 -252
rect 991 -269 995 -256
rect 1015 -257 1019 -245
rect 1050 -249 1054 -237
rect 1044 -253 1054 -249
rect 1019 -261 1024 -257
rect 1087 -261 1090 -257
rect 858 -273 995 -269
rect 858 -278 862 -273
rect 809 -285 811 -281
rect 852 -282 865 -278
rect 809 -293 811 -289
rect 823 -290 832 -286
rect 809 -301 811 -297
rect 823 -302 827 -290
rect 858 -294 862 -282
rect 852 -298 862 -294
rect 827 -306 832 -302
rect 895 -306 898 -302
rect 872 -481 998 -477
rect 872 -486 876 -481
rect 823 -493 825 -489
rect 837 -490 846 -486
rect 872 -490 879 -486
rect 823 -501 825 -497
rect 837 -502 841 -490
rect 872 -494 876 -490
rect 866 -498 876 -494
rect 841 -506 846 -502
rect 899 -506 902 -502
rect 866 -542 976 -538
rect 866 -552 870 -542
rect 817 -559 819 -555
rect 860 -556 873 -552
rect 817 -567 819 -563
rect 831 -564 840 -560
rect 817 -575 819 -571
rect 831 -576 835 -564
rect 866 -568 870 -556
rect 860 -572 870 -568
rect 972 -575 976 -542
rect 994 -567 998 -481
rect 1059 -564 1063 -554
rect 994 -571 1012 -567
rect 1024 -568 1033 -564
rect 1059 -568 1066 -564
rect 835 -580 840 -576
rect 903 -580 906 -576
rect 972 -579 1012 -575
rect 1024 -580 1028 -568
rect 1059 -572 1063 -568
rect 1053 -576 1063 -572
rect 972 -587 1012 -583
rect 1024 -584 1033 -580
rect 972 -604 976 -587
rect 994 -595 1012 -591
rect 994 -624 998 -595
rect 1024 -596 1028 -584
rect 1059 -588 1063 -576
rect 1053 -592 1063 -588
rect 1028 -600 1033 -596
rect 1106 -600 1109 -596
rect 866 -628 998 -624
rect 866 -634 870 -628
rect 817 -641 819 -637
rect 831 -638 840 -634
rect 866 -638 873 -634
rect 817 -649 819 -645
rect 831 -650 835 -638
rect 866 -642 870 -638
rect 860 -646 870 -642
rect 817 -657 819 -653
rect 831 -654 840 -650
rect 817 -665 819 -661
rect 831 -666 835 -654
rect 866 -658 870 -646
rect 860 -662 870 -658
rect 835 -670 840 -666
rect 913 -670 916 -666
rect 874 -895 1023 -891
rect 874 -900 878 -895
rect 825 -907 827 -903
rect 839 -904 848 -900
rect 874 -904 881 -900
rect 825 -915 827 -911
rect 839 -916 843 -904
rect 874 -908 878 -904
rect 868 -912 878 -908
rect 843 -920 848 -916
rect 901 -920 904 -916
rect 868 -952 993 -948
rect 868 -966 872 -952
rect 819 -973 821 -969
rect 862 -970 875 -966
rect 819 -981 821 -977
rect 833 -978 842 -974
rect 819 -989 821 -985
rect 833 -990 837 -978
rect 868 -982 872 -970
rect 862 -986 872 -982
rect 837 -994 842 -990
rect 905 -994 908 -990
rect 959 -1025 971 -1021
rect 868 -1042 946 -1038
rect 868 -1048 872 -1042
rect 942 -1047 946 -1042
rect 967 -1039 971 -1025
rect 989 -1031 993 -952
rect 1019 -1023 1023 -895
rect 1084 -1019 1088 -1010
rect 1078 -1023 1091 -1019
rect 1019 -1027 1037 -1023
rect 1051 -1031 1064 -1027
rect 989 -1035 1037 -1031
rect 967 -1043 1037 -1039
rect 1051 -1043 1055 -1031
rect 1084 -1035 1088 -1023
rect 1078 -1039 1088 -1035
rect 1051 -1047 1064 -1043
rect 819 -1055 821 -1051
rect 833 -1052 842 -1048
rect 868 -1052 875 -1048
rect 942 -1051 1037 -1047
rect 819 -1063 821 -1059
rect 833 -1064 837 -1052
rect 868 -1056 872 -1052
rect 862 -1060 872 -1056
rect 1003 -1059 1037 -1055
rect 1051 -1059 1055 -1047
rect 1084 -1051 1088 -1039
rect 1078 -1055 1088 -1051
rect 819 -1071 821 -1067
rect 833 -1068 842 -1064
rect 819 -1079 821 -1075
rect 833 -1080 837 -1068
rect 868 -1072 872 -1060
rect 862 -1076 872 -1072
rect 837 -1084 842 -1080
rect 915 -1084 918 -1080
rect 1003 -1116 1007 -1059
rect 1055 -1063 1064 -1059
rect 1141 -1063 1144 -1059
rect 869 -1120 1007 -1116
rect 869 -1135 873 -1120
rect 863 -1139 876 -1135
rect 820 -1143 822 -1139
rect 836 -1147 849 -1143
rect 820 -1151 822 -1147
rect 820 -1159 822 -1155
rect 836 -1159 840 -1147
rect 869 -1151 873 -1139
rect 863 -1155 873 -1151
rect 836 -1163 849 -1159
rect 820 -1167 822 -1163
rect 820 -1177 822 -1172
rect 836 -1175 840 -1163
rect 869 -1167 873 -1155
rect 863 -1171 873 -1167
rect 840 -1179 849 -1175
rect 926 -1179 929 -1175
rect 873 -1395 877 -1386
rect 824 -1402 826 -1398
rect 838 -1399 847 -1395
rect 873 -1399 880 -1395
rect 824 -1410 826 -1406
rect 838 -1411 842 -1399
rect 873 -1403 877 -1399
rect 867 -1407 877 -1403
rect 842 -1415 847 -1411
rect 900 -1415 903 -1411
rect 867 -1461 871 -1452
rect 818 -1468 820 -1464
rect 861 -1465 874 -1461
rect 818 -1476 820 -1472
rect 832 -1473 841 -1469
rect 818 -1484 820 -1480
rect 832 -1485 836 -1473
rect 867 -1477 871 -1465
rect 861 -1481 871 -1477
rect 836 -1489 841 -1485
rect 904 -1489 907 -1485
rect 1091 -1527 1095 -1517
rect 867 -1543 871 -1533
rect 1042 -1534 1044 -1530
rect 1056 -1531 1065 -1527
rect 1091 -1531 1098 -1527
rect 1042 -1542 1044 -1538
rect 1056 -1543 1060 -1531
rect 1091 -1535 1095 -1531
rect 1085 -1539 1095 -1535
rect 818 -1550 820 -1546
rect 832 -1547 841 -1543
rect 867 -1547 874 -1543
rect 818 -1558 820 -1554
rect 832 -1559 836 -1547
rect 867 -1551 871 -1547
rect 1042 -1550 1044 -1546
rect 1056 -1547 1065 -1543
rect 861 -1555 871 -1551
rect 818 -1566 820 -1562
rect 832 -1563 841 -1559
rect 818 -1574 820 -1570
rect 832 -1575 836 -1563
rect 867 -1567 871 -1555
rect 1042 -1558 1044 -1554
rect 1056 -1559 1060 -1547
rect 1091 -1551 1095 -1539
rect 1085 -1555 1095 -1551
rect 1042 -1566 1044 -1562
rect 1056 -1563 1065 -1559
rect 861 -1571 871 -1567
rect 1042 -1574 1044 -1570
rect 1056 -1575 1060 -1563
rect 1091 -1567 1095 -1555
rect 1085 -1571 1095 -1567
rect 836 -1579 841 -1575
rect 914 -1579 917 -1575
rect 1060 -1579 1065 -1575
rect 1158 -1579 1161 -1575
rect 868 -1630 872 -1621
rect 862 -1634 875 -1630
rect 819 -1638 821 -1634
rect 835 -1642 848 -1638
rect 819 -1646 821 -1642
rect 819 -1654 821 -1650
rect 835 -1654 839 -1642
rect 868 -1646 872 -1634
rect 862 -1650 872 -1646
rect 835 -1658 848 -1654
rect 819 -1662 821 -1658
rect 819 -1671 821 -1667
rect 835 -1670 839 -1658
rect 868 -1662 872 -1650
rect 862 -1666 872 -1662
rect 839 -1674 848 -1670
rect 925 -1674 928 -1670
rect 864 -1734 868 -1724
rect 815 -1741 817 -1737
rect 829 -1738 838 -1734
rect 864 -1738 871 -1734
rect 815 -1749 817 -1745
rect 829 -1750 833 -1738
rect 864 -1742 868 -1738
rect 858 -1746 868 -1742
rect 815 -1757 817 -1753
rect 829 -1754 838 -1750
rect 815 -1765 817 -1761
rect 829 -1766 833 -1754
rect 864 -1758 868 -1746
rect 858 -1762 868 -1758
rect 829 -1770 838 -1766
rect 815 -1774 817 -1770
rect 815 -1783 817 -1779
rect 829 -1782 833 -1770
rect 864 -1774 868 -1762
rect 858 -1778 868 -1774
rect 833 -1786 838 -1782
rect 931 -1786 934 -1782
rect 0 -2058 155 -2053
<< m2contact >>
rect 219 63 226 70
rect 206 30 211 35
rect 275 41 280 46
rect 342 -48 347 -43
rect 168 -82 173 -77
rect 222 -78 227 -73
rect 325 -89 330 -84
rect 356 -85 361 -80
rect 218 -223 225 -216
rect 209 -244 214 -239
rect 275 -242 280 -237
rect 398 6 403 11
rect 406 -85 411 -80
rect 414 -94 419 -89
rect 218 -361 225 -355
rect 175 -368 180 -363
rect 328 -377 333 -372
rect 363 -373 368 -368
rect 218 -545 225 -538
rect 207 -573 212 -568
rect 275 -571 280 -566
rect 221 -690 226 -685
rect 170 -715 177 -708
rect 332 -703 337 -698
rect 363 -699 368 -694
rect 218 -1025 223 -1020
rect 208 -1064 213 -1059
rect 273 -1060 278 -1055
rect 173 -1187 178 -1182
rect 331 -1188 336 -1183
rect 362 -1184 367 -1179
rect 217 -1522 223 -1516
rect 196 -1554 201 -1549
rect 272 -1550 277 -1545
rect 217 -1669 222 -1664
rect 176 -1677 181 -1672
rect 331 -1674 336 -1669
rect 357 -1674 362 -1669
rect 160 -2024 165 -2019
rect 390 -2024 395 -2019
rect 422 -276 427 -271
rect 430 -373 435 -368
rect 438 -384 443 -379
rect 446 -605 451 -600
rect 454 -699 459 -694
rect 462 -709 467 -704
rect 470 -1061 475 -1056
rect 478 -1184 483 -1179
rect 486 -1247 491 -1242
rect 494 -1585 499 -1580
rect 502 -1679 507 -1674
rect 510 -1738 515 -1733
rect 832 23 837 29
rect 928 -74 933 -68
rect 829 -238 834 -232
rect 1010 -263 1015 -257
rect 829 -312 834 -306
rect 837 -512 842 -506
rect 831 -586 836 -580
rect 1019 -602 1024 -596
rect 831 -676 836 -670
rect 839 -925 844 -920
rect 833 -999 838 -994
rect 833 -1089 838 -1084
rect 1046 -1065 1051 -1059
rect 836 -1185 841 -1179
rect 838 -1421 843 -1415
rect 832 -1495 837 -1489
rect 832 -1585 837 -1579
rect 1051 -1581 1056 -1575
rect 835 -1680 840 -1674
rect 829 -1792 834 -1786
<< pm12contact >>
rect 25 70 30 75
rect 45 70 50 75
rect 117 10 122 15
rect 23 -68 28 -63
rect 43 -68 48 -63
rect 115 -128 120 -123
rect 23 -209 28 -204
rect 43 -209 48 -204
rect 115 -269 120 -264
rect 23 -351 28 -346
rect 43 -351 48 -346
rect 115 -411 120 -406
rect 23 -538 28 -533
rect 43 -538 48 -533
rect 115 -598 120 -593
rect 23 -680 28 -675
rect 43 -680 48 -675
rect 115 -740 120 -735
rect 23 -1028 28 -1023
rect 43 -1028 48 -1023
rect 115 -1088 120 -1083
rect 21 -1169 26 -1164
rect 41 -1169 46 -1164
rect 113 -1229 118 -1224
rect 21 -1518 26 -1513
rect 41 -1518 46 -1513
rect 113 -1578 118 -1573
rect 21 -1659 26 -1654
rect 41 -1659 46 -1654
rect 113 -1719 118 -1714
rect 21 -1988 26 -1983
rect 41 -1988 46 -1983
rect 113 -2048 118 -2043
<< metal2 >>
rect 0 80 28 83
rect 0 48 3 80
rect 24 77 28 80
rect 24 75 50 77
rect 24 74 25 75
rect 30 74 45 75
rect -28 42 3 48
rect 177 63 219 68
rect -28 -78 -22 42
rect 0 12 3 42
rect 0 10 117 12
rect 0 9 121 10
rect -2 -58 26 -55
rect -2 -78 1 -58
rect 22 -61 26 -58
rect 22 -63 48 -61
rect 22 -64 23 -63
rect 28 -64 43 -63
rect 177 -72 182 63
rect -28 -84 1 -78
rect 168 -77 182 -72
rect 206 -73 211 30
rect 275 10 279 41
rect 776 23 832 28
rect 275 6 398 10
rect 776 -43 780 23
rect 347 -48 780 -43
rect 776 -69 780 -48
rect 776 -72 928 -69
rect 206 -78 222 -73
rect -28 -244 -22 -84
rect -2 -126 1 -84
rect 361 -84 406 -80
rect 325 -111 330 -89
rect 358 -94 414 -89
rect 358 -111 363 -94
rect 325 -116 363 -111
rect -2 -128 115 -126
rect -2 -129 119 -128
rect -2 -199 26 -196
rect -2 -244 1 -199
rect 22 -202 26 -199
rect 22 -204 48 -202
rect 22 -205 23 -204
rect 28 -205 43 -204
rect 175 -221 218 -216
rect -28 -250 1 -244
rect -28 -373 -22 -250
rect -2 -267 1 -250
rect -2 -269 115 -267
rect -2 -270 119 -269
rect -2 -341 26 -338
rect -2 -373 1 -341
rect 22 -344 26 -341
rect 22 -346 48 -344
rect 22 -347 23 -346
rect 28 -347 43 -346
rect 175 -363 180 -221
rect 776 -233 780 -72
rect 776 -238 829 -233
rect 209 -261 213 -244
rect 205 -265 213 -261
rect 205 -357 209 -265
rect 275 -272 279 -242
rect 275 -276 422 -272
rect 776 -307 780 -238
rect 1001 -262 1010 -257
rect 776 -312 829 -307
rect 205 -361 218 -357
rect -28 -379 1 -373
rect 368 -373 430 -368
rect -28 -565 -22 -379
rect -2 -409 1 -379
rect -2 -411 115 -409
rect -2 -412 119 -411
rect 328 -424 333 -377
rect 776 -377 780 -312
rect 1001 -377 1006 -262
rect 363 -384 438 -379
rect 776 -382 1006 -377
rect 363 -424 368 -384
rect 328 -429 368 -424
rect 776 -509 780 -382
rect 776 -512 837 -509
rect -2 -528 26 -525
rect -2 -565 1 -528
rect 22 -531 26 -528
rect 22 -533 48 -531
rect 22 -534 23 -533
rect 28 -534 43 -533
rect 170 -545 218 -540
rect -28 -571 1 -565
rect -28 -699 -22 -571
rect -2 -596 1 -571
rect -2 -598 115 -596
rect -2 -599 119 -598
rect -2 -670 26 -667
rect -2 -699 1 -670
rect 22 -673 26 -670
rect 22 -675 48 -673
rect 22 -676 23 -675
rect 28 -676 43 -675
rect -28 -705 1 -699
rect -28 -931 -22 -705
rect -2 -738 1 -705
rect 170 -703 175 -545
rect 207 -577 212 -573
rect 207 -686 211 -577
rect 275 -600 280 -571
rect 776 -583 780 -512
rect 776 -586 831 -583
rect 275 -605 446 -600
rect 776 -673 780 -586
rect 1010 -601 1019 -596
rect 776 -676 831 -673
rect 207 -690 221 -686
rect 170 -708 177 -703
rect 368 -699 454 -694
rect -2 -740 115 -738
rect -2 -741 119 -740
rect 332 -756 337 -703
rect 361 -709 462 -704
rect 361 -756 366 -709
rect 332 -761 366 -756
rect 776 -756 780 -676
rect 1010 -756 1014 -601
rect 776 -761 1014 -756
rect 776 -922 780 -761
rect 776 -925 839 -922
rect -42 -936 -22 -931
rect -28 -1045 -22 -936
rect 776 -996 780 -925
rect 776 -999 833 -996
rect -2 -1018 26 -1015
rect -2 -1045 1 -1018
rect 22 -1021 26 -1018
rect 22 -1023 48 -1021
rect 22 -1024 23 -1023
rect 28 -1024 43 -1023
rect 173 -1025 218 -1020
rect -28 -1051 1 -1045
rect -28 -1199 -22 -1051
rect -2 -1086 1 -1051
rect -2 -1088 115 -1086
rect -2 -1089 119 -1088
rect -4 -1159 24 -1156
rect -4 -1199 -1 -1159
rect 20 -1162 24 -1159
rect 20 -1164 46 -1162
rect 20 -1165 21 -1164
rect 26 -1165 41 -1164
rect 173 -1182 178 -1025
rect 208 -1067 213 -1064
rect 209 -1176 212 -1067
rect 273 -1090 278 -1060
rect 301 -1061 470 -1056
rect 301 -1090 306 -1061
rect 273 -1095 306 -1090
rect 776 -1086 780 -999
rect 1034 -1064 1046 -1060
rect 776 -1089 833 -1086
rect 209 -1179 218 -1176
rect 367 -1184 478 -1179
rect 776 -1182 780 -1089
rect -28 -1205 0 -1199
rect -28 -1555 -22 -1205
rect -4 -1227 -1 -1205
rect -4 -1229 113 -1227
rect -4 -1230 117 -1229
rect 331 -1242 336 -1188
rect 776 -1185 836 -1182
rect 331 -1247 486 -1242
rect 776 -1260 780 -1185
rect 1034 -1260 1038 -1064
rect 776 -1264 1038 -1260
rect 776 -1417 780 -1264
rect 776 -1421 838 -1417
rect 776 -1492 780 -1421
rect 776 -1495 832 -1492
rect -4 -1508 24 -1505
rect -4 -1555 -1 -1508
rect 20 -1511 24 -1508
rect 20 -1513 46 -1511
rect 20 -1514 21 -1513
rect 26 -1514 41 -1513
rect 177 -1520 217 -1516
rect -28 -1561 0 -1555
rect -28 -1686 -22 -1561
rect -4 -1576 -1 -1561
rect -4 -1578 113 -1576
rect -4 -1579 117 -1578
rect -4 -1649 24 -1646
rect -4 -1686 -1 -1649
rect 20 -1652 24 -1649
rect 20 -1654 46 -1652
rect 20 -1655 21 -1654
rect 26 -1655 41 -1654
rect 177 -1668 181 -1520
rect 176 -1672 181 -1668
rect 196 -1664 201 -1554
rect 272 -1580 277 -1550
rect 272 -1585 494 -1580
rect 776 -1582 780 -1495
rect 776 -1585 832 -1582
rect 1041 -1580 1051 -1576
rect 196 -1669 217 -1664
rect -28 -1692 0 -1686
rect -28 -2009 -22 -1692
rect -4 -1717 -1 -1692
rect -4 -1719 113 -1717
rect -4 -1720 117 -1719
rect 331 -1733 336 -1674
rect 357 -1679 502 -1674
rect 776 -1677 780 -1585
rect 776 -1680 835 -1677
rect 331 -1738 510 -1733
rect 776 -1789 780 -1680
rect 776 -1792 829 -1789
rect 776 -1876 780 -1792
rect 1041 -1876 1045 -1580
rect 776 -1880 1045 -1876
rect -4 -1978 24 -1975
rect -4 -2009 -1 -1978
rect 20 -1981 24 -1978
rect 20 -1983 46 -1981
rect 20 -1984 21 -1983
rect 26 -1984 41 -1983
rect -28 -2015 0 -2009
rect -4 -2046 -1 -2015
rect 165 -2024 390 -2019
rect -4 -2048 113 -2046
rect -4 -2049 117 -2048
<< m3contact >>
rect 83 -1511 88 -1506
<< m123contact >>
rect 162 90 167 95
rect 45 82 50 87
rect 87 80 92 85
rect 28 38 33 43
rect 160 -48 165 -43
rect 43 -56 48 -51
rect 85 -61 90 -56
rect 232 54 237 59
rect 399 43 404 48
rect 814 43 819 48
rect 391 32 396 37
rect 814 32 819 37
rect 894 24 899 29
rect 523 11 528 16
rect 333 -50 338 -45
rect 415 -64 420 -59
rect 909 -64 914 -59
rect 523 -78 528 -73
rect 234 -92 239 -87
rect 26 -100 31 -95
rect 160 -189 165 -184
rect 43 -197 48 -192
rect 85 -202 90 -197
rect 26 -241 31 -236
rect 160 -331 165 -326
rect 43 -339 48 -334
rect 85 -344 90 -339
rect 423 -218 428 -213
rect 232 -229 237 -224
rect 407 -229 412 -224
rect 990 -73 995 -68
rect 810 -218 815 -213
rect 810 -229 815 -224
rect 891 -237 896 -232
rect 523 -247 528 -242
rect 439 -263 444 -257
rect 423 -285 428 -280
rect 399 -293 404 -288
rect 391 -302 396 -297
rect 981 -248 987 -242
rect 804 -284 809 -279
rect 804 -293 809 -288
rect 804 -302 809 -297
rect 895 -311 900 -306
rect 523 -321 528 -316
rect 336 -337 341 -332
rect 234 -375 239 -370
rect 26 -383 31 -378
rect 1087 -266 1092 -261
rect 447 -494 452 -489
rect 431 -504 436 -499
rect 818 -493 823 -488
rect 818 -503 823 -498
rect 899 -511 904 -506
rect 160 -518 165 -513
rect 43 -526 48 -521
rect 523 -525 528 -520
rect 85 -531 90 -526
rect 26 -570 31 -565
rect 160 -660 165 -655
rect 43 -668 48 -663
rect 85 -673 90 -668
rect 232 -558 237 -553
rect 447 -559 452 -554
rect 423 -568 428 -563
rect 407 -577 412 -572
rect 812 -558 817 -553
rect 812 -567 817 -562
rect 812 -576 817 -571
rect 903 -585 908 -580
rect 523 -595 528 -590
rect 463 -609 468 -604
rect 447 -641 452 -636
rect 423 -650 428 -645
rect 399 -659 404 -654
rect 336 -664 341 -659
rect 391 -668 396 -663
rect 971 -610 977 -604
rect 812 -640 817 -635
rect 812 -649 817 -644
rect 812 -658 817 -653
rect 812 -667 817 -662
rect 913 -675 918 -670
rect 523 -685 528 -680
rect 26 -712 31 -707
rect 234 -704 239 -699
rect 1106 -605 1111 -600
rect 471 -907 476 -902
rect 455 -916 460 -911
rect 820 -906 825 -901
rect 820 -915 825 -910
rect 901 -925 906 -920
rect 523 -930 528 -925
rect 471 -973 476 -968
rect 447 -982 452 -977
rect 431 -991 436 -985
rect 814 -972 819 -967
rect 814 -981 819 -976
rect 814 -990 819 -985
rect 905 -999 910 -994
rect 160 -1008 165 -1003
rect 523 -1009 528 -1004
rect 43 -1016 48 -1011
rect 85 -1021 90 -1016
rect 26 -1060 31 -1055
rect 158 -1149 163 -1144
rect 41 -1157 46 -1152
rect 83 -1162 88 -1157
rect 487 -1026 492 -1020
rect 471 -1038 476 -1032
rect 232 -1047 237 -1042
rect 447 -1050 452 -1045
rect 423 -1073 428 -1067
rect 407 -1082 412 -1077
rect 954 -1026 959 -1020
rect 814 -1054 819 -1049
rect 814 -1063 819 -1058
rect 814 -1072 819 -1067
rect 814 -1081 819 -1076
rect 915 -1089 920 -1084
rect 523 -1099 528 -1094
rect 471 -1143 476 -1138
rect 335 -1149 340 -1144
rect 447 -1152 452 -1147
rect 390 -1158 395 -1152
rect 423 -1161 428 -1156
rect 399 -1170 404 -1165
rect 815 -1142 820 -1137
rect 815 -1151 820 -1146
rect 815 -1160 820 -1155
rect 815 -1169 820 -1164
rect 815 -1178 820 -1173
rect 232 -1193 237 -1188
rect 24 -1201 29 -1196
rect 926 -1184 931 -1179
rect 523 -1194 528 -1189
rect 1141 -1068 1146 -1063
rect 495 -1403 500 -1398
rect 479 -1412 484 -1407
rect 819 -1402 824 -1397
rect 819 -1411 824 -1406
rect 900 -1420 905 -1415
rect 523 -1430 528 -1425
rect 495 -1468 500 -1463
rect 471 -1477 476 -1472
rect 455 -1486 460 -1481
rect 813 -1467 818 -1462
rect 813 -1476 818 -1471
rect 813 -1485 818 -1480
rect 158 -1498 163 -1493
rect 904 -1494 909 -1489
rect 41 -1506 46 -1501
rect 523 -1504 528 -1499
rect 24 -1550 29 -1545
rect 158 -1639 163 -1634
rect 41 -1647 46 -1642
rect 83 -1652 88 -1647
rect 232 -1537 237 -1532
rect 495 -1550 500 -1545
rect 471 -1559 476 -1554
rect 447 -1568 452 -1563
rect 430 -1573 436 -1568
rect 813 -1549 818 -1544
rect 813 -1558 818 -1553
rect 813 -1567 818 -1562
rect 813 -1576 818 -1571
rect 914 -1584 919 -1579
rect 523 -1594 528 -1589
rect 335 -1635 340 -1630
rect 495 -1638 500 -1633
rect 471 -1647 476 -1642
rect 447 -1656 452 -1651
rect 407 -1664 412 -1658
rect 423 -1665 428 -1660
rect 231 -1683 236 -1678
rect 24 -1691 29 -1686
rect 814 -1637 819 -1632
rect 814 -1646 819 -1641
rect 814 -1655 819 -1650
rect 814 -1664 819 -1659
rect 814 -1673 819 -1668
rect 925 -1679 930 -1674
rect 523 -1689 528 -1684
rect 495 -1747 500 -1742
rect 471 -1756 476 -1751
rect 447 -1765 452 -1760
rect 399 -1775 404 -1770
rect 423 -1774 428 -1769
rect 391 -1791 396 -1786
rect 810 -1740 815 -1735
rect 810 -1749 815 -1744
rect 810 -1758 815 -1753
rect 810 -1767 815 -1762
rect 810 -1776 815 -1771
rect 810 -1785 815 -1780
rect 931 -1791 936 -1786
rect 523 -1801 528 -1796
rect 1158 -1584 1163 -1579
rect 158 -1968 163 -1963
rect 41 -1976 46 -1971
rect 83 -1981 88 -1976
rect 24 -2020 29 -2015
<< metal3 >>
rect 167 90 190 94
rect 35 82 45 87
rect 35 43 38 82
rect 75 80 87 83
rect 33 38 39 43
rect 33 -56 43 -51
rect 33 -95 36 -56
rect 75 -58 78 80
rect 186 59 190 90
rect 186 54 232 59
rect 186 -44 190 54
rect 404 43 814 46
rect 396 32 814 35
rect 894 15 898 24
rect 528 11 898 15
rect 165 -45 190 -44
rect 165 -48 333 -45
rect 186 -49 333 -48
rect 75 -61 85 -58
rect 31 -100 37 -95
rect 33 -197 43 -192
rect 33 -236 36 -197
rect 75 -199 78 -61
rect 186 -87 190 -49
rect 420 -64 909 -61
rect 528 -78 995 -73
rect 186 -92 234 -87
rect 186 -185 190 -92
rect 165 -189 190 -185
rect 75 -202 85 -199
rect 31 -241 37 -236
rect 33 -339 43 -334
rect 33 -378 36 -339
rect 75 -341 78 -202
rect 186 -224 190 -189
rect 428 -218 810 -215
rect 186 -229 232 -224
rect 412 -229 810 -226
rect 186 -327 190 -229
rect 891 -242 896 -237
rect 528 -247 896 -242
rect 957 -248 981 -242
rect 957 -257 963 -248
rect 444 -263 963 -257
rect 428 -284 804 -281
rect 404 -293 804 -290
rect 396 -302 804 -299
rect 895 -316 900 -311
rect 1087 -316 1092 -266
rect 528 -321 1092 -316
rect 165 -331 190 -327
rect 186 -332 190 -331
rect 186 -336 336 -332
rect 75 -344 85 -341
rect 31 -383 37 -378
rect 33 -526 43 -521
rect 33 -565 36 -526
rect 75 -528 78 -344
rect 186 -370 190 -336
rect 186 -375 234 -370
rect 186 -514 190 -375
rect 452 -493 818 -490
rect 436 -503 818 -500
rect 165 -518 190 -514
rect 75 -531 85 -528
rect 31 -570 37 -565
rect 33 -668 43 -663
rect 33 -707 36 -668
rect 75 -670 78 -531
rect 186 -553 190 -518
rect 899 -520 904 -511
rect 528 -525 904 -520
rect 186 -558 232 -553
rect 186 -656 190 -558
rect 452 -558 812 -555
rect 428 -567 812 -564
rect 412 -576 812 -573
rect 903 -590 908 -585
rect 528 -595 908 -590
rect 468 -609 971 -605
rect 452 -640 812 -637
rect 428 -649 812 -646
rect 165 -659 190 -656
rect 404 -658 812 -655
rect 165 -660 336 -659
rect 186 -663 336 -660
rect 75 -673 85 -670
rect 31 -712 37 -707
rect 75 -881 78 -673
rect 186 -699 190 -663
rect 396 -667 812 -664
rect 913 -678 918 -675
rect 1106 -678 1111 -605
rect 913 -680 1111 -678
rect 528 -683 1111 -680
rect 528 -685 918 -683
rect 186 -704 234 -699
rect 186 -840 190 -704
rect 181 -844 190 -840
rect 63 -885 78 -881
rect 33 -1016 43 -1011
rect 33 -1055 36 -1016
rect 75 -1018 78 -885
rect 186 -1004 190 -844
rect 476 -906 820 -903
rect 460 -915 820 -912
rect 528 -930 906 -925
rect 476 -972 814 -969
rect 452 -981 814 -978
rect 436 -990 814 -987
rect 905 -1004 910 -999
rect 165 -1008 190 -1004
rect 75 -1021 85 -1018
rect 31 -1060 37 -1055
rect 31 -1157 41 -1152
rect 31 -1196 34 -1157
rect 75 -1159 78 -1021
rect 186 -1042 190 -1008
rect 528 -1009 910 -1004
rect 492 -1026 954 -1020
rect 476 -1037 529 -1034
rect 186 -1047 232 -1042
rect 186 -1144 190 -1047
rect 452 -1049 518 -1046
rect 515 -1060 518 -1049
rect 526 -1051 529 -1037
rect 526 -1054 814 -1051
rect 515 -1063 814 -1060
rect 428 -1072 814 -1069
rect 412 -1081 814 -1078
rect 915 -1090 920 -1089
rect 1141 -1090 1146 -1068
rect 915 -1094 1146 -1090
rect 528 -1095 1146 -1094
rect 528 -1099 920 -1095
rect 476 -1142 815 -1139
rect 186 -1145 335 -1144
rect 163 -1148 335 -1145
rect 163 -1149 190 -1148
rect 75 -1162 83 -1159
rect 29 -1201 35 -1196
rect 31 -1506 41 -1501
rect 31 -1545 34 -1506
rect 75 -1508 78 -1162
rect 186 -1188 190 -1149
rect 452 -1151 815 -1148
rect 392 -1175 395 -1158
rect 428 -1160 815 -1157
rect 404 -1169 815 -1166
rect 392 -1178 815 -1175
rect 186 -1193 232 -1188
rect 926 -1189 931 -1184
rect 186 -1494 190 -1193
rect 528 -1194 931 -1189
rect 500 -1402 819 -1399
rect 484 -1411 819 -1408
rect 900 -1425 905 -1420
rect 528 -1430 909 -1425
rect 500 -1467 813 -1464
rect 476 -1476 813 -1473
rect 460 -1485 813 -1482
rect 163 -1498 190 -1494
rect 75 -1511 83 -1508
rect 29 -1550 35 -1545
rect 31 -1647 41 -1642
rect 31 -1686 34 -1647
rect 75 -1649 78 -1511
rect 186 -1532 190 -1498
rect 904 -1499 909 -1494
rect 528 -1504 917 -1499
rect 186 -1537 232 -1532
rect 186 -1630 190 -1537
rect 500 -1549 813 -1546
rect 476 -1558 813 -1555
rect 452 -1567 813 -1564
rect 431 -1576 813 -1573
rect 914 -1589 919 -1584
rect 1158 -1589 1163 -1584
rect 528 -1594 1163 -1589
rect 186 -1634 335 -1630
rect 186 -1635 190 -1634
rect 163 -1639 190 -1635
rect 500 -1637 814 -1634
rect 75 -1652 83 -1649
rect 29 -1691 35 -1686
rect 31 -1976 41 -1971
rect 31 -2015 34 -1976
rect 75 -1978 78 -1652
rect 186 -1678 190 -1639
rect 476 -1646 814 -1643
rect 452 -1655 814 -1652
rect 407 -1670 410 -1664
rect 428 -1664 814 -1661
rect 407 -1673 814 -1670
rect 186 -1683 231 -1678
rect 186 -1964 190 -1683
rect 925 -1684 930 -1679
rect 528 -1689 930 -1684
rect 527 -1740 810 -1737
rect 527 -1743 530 -1740
rect 500 -1746 530 -1743
rect 534 -1749 810 -1746
rect 534 -1752 537 -1749
rect 476 -1755 537 -1752
rect 541 -1758 810 -1755
rect 541 -1761 544 -1758
rect 452 -1764 544 -1761
rect 549 -1767 810 -1764
rect 549 -1770 552 -1767
rect 428 -1773 552 -1770
rect 399 -1779 402 -1775
rect 556 -1776 810 -1773
rect 556 -1779 559 -1776
rect 399 -1782 559 -1779
rect 565 -1785 810 -1782
rect 565 -1787 568 -1785
rect 396 -1790 568 -1787
rect 931 -1796 936 -1791
rect 528 -1801 936 -1796
rect 163 -1968 190 -1964
rect 75 -1981 83 -1978
rect 29 -2020 35 -2015
<< metal4 >>
rect 437 29 441 33
<< labels >>
rlabel metal1 17 74 21 77 1 a0
rlabel metal1 15 -64 19 -61 1 b0
rlabel metal1 15 -205 19 -202 1 a1
rlabel metal1 15 -347 19 -344 1 b1
rlabel metal1 15 -534 19 -531 1 a2
rlabel metal1 15 -676 19 -673 1 b2
rlabel metal1 15 -1024 19 -1021 1 a3
rlabel metal1 13 -1165 17 -1162 1 b3
rlabel metal1 13 -1514 17 -1511 1 a4
rlabel metal1 13 -1655 17 -1652 1 b4
rlabel metal1 13 -1984 17 -1981 1 c0
rlabel metal2 -42 -936 -28 -931 1 clk
rlabel metal3 63 -885 75 -881 1 rst
rlabel metal1 -9 -1382 -4 -1378 1 gnd
rlabel metal3 181 -844 186 -840 1 vdd
rlabel metal1 135 35 138 39 1 qb0
rlabel metal1 159 35 162 39 1 q0
rlabel metal1 136 -103 139 -99 1 qb5
rlabel metal1 158 -103 161 -99 1 q5
rlabel metal1 138 -244 141 -240 1 qb1
rlabel metal1 158 -244 161 -240 1 q1
rlabel metal1 133 -386 136 -382 1 qb6
rlabel metal1 158 -386 161 -382 1 q6
rlabel metal1 134 -573 137 -569 1 qb2
rlabel metal1 157 -573 160 -569 1 q2
rlabel metal1 134 -715 137 -711 1 qb7
rlabel metal1 157 -715 160 -711 1 q7
rlabel metal1 135 -1063 138 -1059 1 qb3
rlabel metal1 157 -1063 160 -1059 1 q3
rlabel metal1 133 -1204 136 -1200 1 qb8
rlabel metal1 155 -1204 158 -1200 1 q8
rlabel metal1 135 -1553 138 -1549 1 qb4
rlabel metal1 155 -1553 158 -1549 1 q4
rlabel metal1 134 -1694 137 -1690 1 qb9
rlabel metal1 155 -1694 158 -1690 1 q9
rlabel metal1 155 -2023 158 -2019 1 qc0
rlabel metal1 132 -2023 135 -2019 1 qbc0
rlabel metal1 275 46 279 50 1 p0
rlabel metal1 325 -84 328 -80 1 g0_bar
rlabel metal1 353 -84 356 -80 1 g0
rlabel metal1 275 -237 278 -233 1 p1
rlabel metal1 329 -372 332 -368 1 g1_bar
rlabel metal1 359 -372 362 -368 1 g1
rlabel metal1 275 -566 278 -562 1 p2
rlabel metal1 335 -698 338 -694 1 g2_bar
rlabel metal1 355 -698 358 -694 1 g2
rlabel metal1 273 -1055 276 -1051 1 p3
rlabel metal1 334 -1183 337 -1179 1 g3_bar
rlabel metal1 356 -1183 359 -1179 1 g3
rlabel metal1 272 -1545 275 -1541 1 p4
rlabel metal1 334 -1669 337 -1665 1 g4_bar
rlabel metal1 359 -1669 362 -1665 1 g4
rlabel metal1 963 -42 967 -39 1 c1
rlabel metal1 1050 -227 1054 -224 1 c2
rlabel metal1 1059 -557 1063 -554 1 c3
rlabel metal1 1084 -1012 1088 -1010 1 c4
rlabel metal1 1091 -1519 1095 -1517 1 cout
<< end >>
