magic
tech scmos
timestamp 1763385314
<< nwell >>
rect 0 0 56 40
<< pdiffusion >>
rect 10 6 50 20
<< pdcontact >>
rect 6 6 10 20
<< end >>
