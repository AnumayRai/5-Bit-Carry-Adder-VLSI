magic
tech scmos
timestamp 1764698668
<< nwell >>
rect 48 2098 205 2159
rect 305 2155 317 2159
rect 272 2115 368 2155
rect 1189 2137 1201 2141
rect 114 2097 147 2098
rect 272 2078 296 2115
rect 704 2081 744 2113
rect 1156 2097 1252 2137
rect 1156 2060 1180 2097
rect 1469 2049 1626 2110
rect 1535 2048 1568 2049
rect 46 1960 203 2021
rect 276 1961 316 1993
rect 374 1979 398 2016
rect 800 1984 840 2016
rect 112 1959 145 1960
rect 46 1819 203 1880
rect 305 1872 317 1876
rect 272 1832 368 1872
rect 112 1818 145 1819
rect 272 1795 296 1832
rect 701 1820 741 1852
rect 1187 1841 1199 1845
rect 887 1791 927 1831
rect 1154 1801 1250 1841
rect 695 1746 735 1786
rect 1154 1764 1178 1801
rect 1469 1787 1626 1848
rect 1535 1786 1568 1787
rect 46 1677 203 1738
rect 276 1678 316 1710
rect 377 1691 401 1728
rect 112 1676 145 1677
rect 46 1490 203 1551
rect 305 1543 317 1547
rect 709 1546 749 1578
rect 272 1503 368 1543
rect 112 1489 145 1490
rect 272 1466 296 1503
rect 703 1472 743 1512
rect 896 1452 936 1500
rect 1187 1481 1199 1485
rect 1154 1441 1250 1481
rect 46 1348 203 1409
rect 276 1349 316 1381
rect 377 1365 401 1402
rect 703 1382 743 1430
rect 1154 1404 1178 1441
rect 1469 1420 1626 1481
rect 1535 1419 1568 1420
rect 112 1347 145 1348
rect 711 1132 751 1164
rect 46 1000 203 1061
rect 705 1058 745 1098
rect 1187 1066 1199 1070
rect 303 1054 315 1058
rect 270 1014 366 1054
rect 112 999 145 1000
rect 270 977 294 1014
rect 705 968 745 1016
rect 921 989 961 1045
rect 1154 1026 1250 1066
rect 1154 989 1178 1026
rect 1469 1002 1626 1063
rect 1535 1001 1568 1002
rect 44 859 201 920
rect 274 860 314 892
rect 376 880 400 917
rect 706 873 746 929
rect 110 858 143 859
rect 710 637 750 669
rect 44 510 201 571
rect 302 564 314 568
rect 269 524 365 564
rect 704 563 744 603
rect 110 509 143 510
rect 269 487 293 524
rect 704 473 744 521
rect 928 473 968 537
rect 1187 526 1199 530
rect 1154 486 1250 526
rect 1154 449 1178 486
rect 44 369 201 430
rect 273 370 313 402
rect 376 394 400 431
rect 705 378 745 434
rect 1469 426 1626 487
rect 1535 425 1568 426
rect 110 368 143 369
rect 701 266 741 330
rect 1469 136 1626 197
rect 1535 135 1568 136
rect 44 40 201 101
rect 110 39 143 40
<< ntransistor >>
rect 59 2081 61 2091
rect 89 2081 91 2091
rect 97 2081 99 2091
rect 152 2077 154 2087
rect 160 2077 162 2087
rect 192 2080 194 2090
rect 307 2098 309 2108
rect 330 2092 332 2102
rect 751 2100 771 2102
rect 751 2092 771 2094
rect 283 2060 285 2070
rect 1191 2080 1193 2090
rect 1214 2074 1216 2084
rect 1167 2042 1169 2052
rect 1480 2032 1482 2042
rect 1510 2032 1512 2042
rect 1518 2032 1520 2042
rect 1573 2028 1575 2038
rect 1581 2028 1583 2038
rect 1613 2031 1615 2041
rect 847 2003 867 2005
rect 847 1995 867 1997
rect 323 1980 343 1982
rect 323 1972 343 1974
rect 57 1943 59 1953
rect 87 1943 89 1953
rect 95 1943 97 1953
rect 385 1961 387 1971
rect 150 1939 152 1949
rect 158 1939 160 1949
rect 190 1942 192 1952
rect 748 1839 768 1841
rect 748 1831 768 1833
rect 57 1802 59 1812
rect 87 1802 89 1812
rect 95 1802 97 1812
rect 150 1798 152 1808
rect 158 1798 160 1808
rect 190 1801 192 1811
rect 307 1815 309 1825
rect 330 1809 332 1819
rect 934 1818 964 1820
rect 934 1810 964 1812
rect 934 1802 964 1804
rect 283 1777 285 1787
rect 742 1773 772 1775
rect 1189 1784 1191 1794
rect 1212 1778 1214 1788
rect 1480 1770 1482 1780
rect 1510 1770 1512 1780
rect 1518 1770 1520 1780
rect 742 1765 772 1767
rect 742 1757 772 1759
rect 1573 1766 1575 1776
rect 1581 1766 1583 1776
rect 1613 1769 1615 1779
rect 1165 1746 1167 1756
rect 323 1697 343 1699
rect 323 1689 343 1691
rect 57 1660 59 1670
rect 87 1660 89 1670
rect 95 1660 97 1670
rect 388 1673 390 1683
rect 150 1656 152 1666
rect 158 1656 160 1666
rect 190 1659 192 1669
rect 756 1565 776 1567
rect 756 1557 776 1559
rect 750 1499 780 1501
rect 57 1473 59 1483
rect 87 1473 89 1483
rect 95 1473 97 1483
rect 150 1469 152 1479
rect 158 1469 160 1479
rect 190 1472 192 1482
rect 307 1486 309 1496
rect 750 1491 780 1493
rect 330 1480 332 1490
rect 943 1487 983 1489
rect 750 1483 780 1485
rect 943 1479 983 1481
rect 943 1471 983 1473
rect 943 1463 983 1465
rect 283 1448 285 1458
rect 750 1417 790 1419
rect 750 1409 790 1411
rect 1189 1424 1191 1434
rect 1212 1418 1214 1428
rect 750 1401 790 1403
rect 1480 1403 1482 1413
rect 1510 1403 1512 1413
rect 1518 1403 1520 1413
rect 1573 1399 1575 1409
rect 1581 1399 1583 1409
rect 1613 1402 1615 1412
rect 750 1393 790 1395
rect 1165 1386 1167 1396
rect 323 1368 343 1370
rect 323 1360 343 1362
rect 57 1331 59 1341
rect 87 1331 89 1341
rect 95 1331 97 1341
rect 388 1347 390 1357
rect 150 1327 152 1337
rect 158 1327 160 1337
rect 190 1330 192 1340
rect 758 1151 778 1153
rect 758 1143 778 1145
rect 752 1085 782 1087
rect 752 1077 782 1079
rect 752 1069 782 1071
rect 968 1032 1018 1034
rect 968 1024 1018 1026
rect 968 1016 1018 1018
rect 57 983 59 993
rect 87 983 89 993
rect 95 983 97 993
rect 150 979 152 989
rect 158 979 160 989
rect 190 982 192 992
rect 305 997 307 1007
rect 968 1008 1018 1010
rect 752 1003 792 1005
rect 328 991 330 1001
rect 968 1000 1018 1002
rect 752 995 792 997
rect 1189 1009 1191 1019
rect 1212 1003 1214 1013
rect 752 987 792 989
rect 1480 985 1482 995
rect 1510 985 1512 995
rect 1518 985 1520 995
rect 1573 981 1575 991
rect 1581 981 1583 991
rect 1613 984 1615 994
rect 752 979 792 981
rect 1165 971 1167 981
rect 281 959 283 969
rect 753 916 803 918
rect 753 908 803 910
rect 753 900 803 902
rect 753 892 803 894
rect 321 879 341 881
rect 321 871 341 873
rect 753 884 803 886
rect 55 842 57 852
rect 85 842 87 852
rect 93 842 95 852
rect 387 862 389 872
rect 148 838 150 848
rect 156 838 158 848
rect 188 841 190 851
rect 757 656 777 658
rect 757 648 777 650
rect 751 590 781 592
rect 751 582 781 584
rect 751 574 781 576
rect 975 524 1035 526
rect 55 493 57 503
rect 85 493 87 503
rect 93 493 95 503
rect 148 489 150 499
rect 156 489 158 499
rect 188 492 190 502
rect 304 507 306 517
rect 975 516 1035 518
rect 327 501 329 511
rect 751 508 791 510
rect 975 508 1035 510
rect 751 500 791 502
rect 975 500 1035 502
rect 751 492 791 494
rect 975 492 1035 494
rect 751 484 791 486
rect 975 484 1035 486
rect 280 469 282 479
rect 1189 469 1191 479
rect 1212 463 1214 473
rect 1165 431 1167 441
rect 752 421 802 423
rect 752 413 802 415
rect 1480 409 1482 419
rect 1510 409 1512 419
rect 1518 409 1520 419
rect 752 405 802 407
rect 1573 405 1575 415
rect 1581 405 1583 415
rect 1613 408 1615 418
rect 320 389 340 391
rect 752 397 802 399
rect 752 389 802 391
rect 320 381 340 383
rect 387 376 389 386
rect 55 352 57 362
rect 85 352 87 362
rect 93 352 95 362
rect 148 348 150 358
rect 156 348 158 358
rect 188 351 190 361
rect 748 317 808 319
rect 748 309 808 311
rect 748 301 808 303
rect 748 293 808 295
rect 748 285 808 287
rect 748 277 808 279
rect 1480 119 1482 129
rect 1510 119 1512 129
rect 1518 119 1520 129
rect 1573 115 1575 125
rect 1581 115 1583 125
rect 1613 118 1615 128
rect 55 23 57 33
rect 85 23 87 33
rect 93 23 95 33
rect 148 19 150 29
rect 156 19 158 29
rect 188 22 190 32
<< ptransistor >>
rect 59 2104 61 2124
rect 67 2104 69 2124
rect 89 2104 91 2124
rect 97 2104 99 2124
rect 129 2107 131 2127
rect 152 2120 154 2140
rect 192 2104 194 2124
rect 307 2121 309 2141
rect 330 2121 332 2141
rect 283 2084 285 2104
rect 1191 2103 1193 2123
rect 1214 2103 1216 2123
rect 718 2100 738 2102
rect 718 2092 738 2094
rect 1167 2066 1169 2086
rect 1480 2055 1482 2075
rect 1488 2055 1490 2075
rect 1510 2055 1512 2075
rect 1518 2055 1520 2075
rect 1550 2058 1552 2078
rect 1573 2071 1575 2091
rect 1613 2055 1615 2075
rect 57 1966 59 1986
rect 65 1966 67 1986
rect 87 1966 89 1986
rect 95 1966 97 1986
rect 127 1969 129 1989
rect 150 1982 152 2002
rect 190 1966 192 1986
rect 385 1985 387 2005
rect 814 2003 834 2005
rect 814 1995 834 1997
rect 290 1980 310 1982
rect 290 1972 310 1974
rect 57 1825 59 1845
rect 65 1825 67 1845
rect 87 1825 89 1845
rect 95 1825 97 1845
rect 127 1828 129 1848
rect 150 1841 152 1861
rect 190 1825 192 1845
rect 307 1838 309 1858
rect 330 1838 332 1858
rect 715 1839 735 1841
rect 715 1831 735 1833
rect 283 1801 285 1821
rect 901 1818 921 1820
rect 901 1810 921 1812
rect 1189 1807 1191 1827
rect 1212 1807 1214 1827
rect 901 1802 921 1804
rect 709 1773 729 1775
rect 1165 1770 1167 1790
rect 1480 1793 1482 1813
rect 1488 1793 1490 1813
rect 1510 1793 1512 1813
rect 1518 1793 1520 1813
rect 1550 1796 1552 1816
rect 1573 1809 1575 1829
rect 1613 1793 1615 1813
rect 709 1765 729 1767
rect 709 1757 729 1759
rect 57 1683 59 1703
rect 65 1683 67 1703
rect 87 1683 89 1703
rect 95 1683 97 1703
rect 127 1686 129 1706
rect 150 1699 152 1719
rect 190 1683 192 1703
rect 290 1697 310 1699
rect 388 1697 390 1717
rect 290 1689 310 1691
rect 723 1565 743 1567
rect 723 1557 743 1559
rect 57 1496 59 1516
rect 65 1496 67 1516
rect 87 1496 89 1516
rect 95 1496 97 1516
rect 127 1499 129 1519
rect 150 1512 152 1532
rect 190 1496 192 1516
rect 307 1509 309 1529
rect 330 1509 332 1529
rect 717 1499 737 1501
rect 283 1472 285 1492
rect 717 1491 737 1493
rect 910 1487 930 1489
rect 717 1483 737 1485
rect 910 1479 930 1481
rect 910 1471 930 1473
rect 910 1463 930 1465
rect 1189 1447 1191 1467
rect 1212 1447 1214 1467
rect 717 1417 737 1419
rect 717 1409 737 1411
rect 1165 1410 1167 1430
rect 1480 1426 1482 1446
rect 1488 1426 1490 1446
rect 1510 1426 1512 1446
rect 1518 1426 1520 1446
rect 1550 1429 1552 1449
rect 1573 1442 1575 1462
rect 1613 1426 1615 1446
rect 717 1401 737 1403
rect 717 1393 737 1395
rect 57 1354 59 1374
rect 65 1354 67 1374
rect 87 1354 89 1374
rect 95 1354 97 1374
rect 127 1357 129 1377
rect 150 1370 152 1390
rect 190 1354 192 1374
rect 388 1371 390 1391
rect 290 1368 310 1370
rect 290 1360 310 1362
rect 725 1151 745 1153
rect 725 1143 745 1145
rect 719 1085 739 1087
rect 719 1077 739 1079
rect 719 1069 739 1071
rect 57 1006 59 1026
rect 65 1006 67 1026
rect 87 1006 89 1026
rect 95 1006 97 1026
rect 127 1009 129 1029
rect 150 1022 152 1042
rect 190 1006 192 1026
rect 305 1020 307 1040
rect 328 1020 330 1040
rect 941 1032 955 1034
rect 1189 1032 1191 1052
rect 1212 1032 1214 1052
rect 941 1024 955 1026
rect 941 1016 955 1018
rect 281 983 283 1003
rect 941 1008 955 1010
rect 719 1003 739 1005
rect 941 1000 955 1002
rect 719 995 739 997
rect 1165 995 1167 1015
rect 1480 1008 1482 1028
rect 1488 1008 1490 1028
rect 1510 1008 1512 1028
rect 1518 1008 1520 1028
rect 1550 1011 1552 1031
rect 1573 1024 1575 1044
rect 1613 1008 1615 1028
rect 719 987 739 989
rect 719 979 739 981
rect 726 916 740 918
rect 726 908 740 910
rect 55 865 57 885
rect 63 865 65 885
rect 85 865 87 885
rect 93 865 95 885
rect 125 868 127 888
rect 148 881 150 901
rect 387 886 389 906
rect 726 900 740 902
rect 726 892 740 894
rect 188 865 190 885
rect 288 879 308 881
rect 288 871 308 873
rect 726 884 740 886
rect 724 656 744 658
rect 724 648 744 650
rect 718 590 738 592
rect 718 582 738 584
rect 718 574 738 576
rect 55 516 57 536
rect 63 516 65 536
rect 85 516 87 536
rect 93 516 95 536
rect 125 519 127 539
rect 148 532 150 552
rect 188 516 190 536
rect 304 530 306 550
rect 327 530 329 550
rect 942 524 962 526
rect 280 493 282 513
rect 942 516 962 518
rect 718 508 738 510
rect 942 508 962 510
rect 718 500 738 502
rect 942 500 962 502
rect 718 492 738 494
rect 942 492 962 494
rect 1189 492 1191 512
rect 1212 492 1214 512
rect 718 484 738 486
rect 942 484 962 486
rect 1165 455 1167 475
rect 1480 432 1482 452
rect 1488 432 1490 452
rect 1510 432 1512 452
rect 1518 432 1520 452
rect 1550 435 1552 455
rect 1573 448 1575 468
rect 725 421 739 423
rect 55 375 57 395
rect 63 375 65 395
rect 85 375 87 395
rect 93 375 95 395
rect 125 378 127 398
rect 148 391 150 411
rect 387 400 389 420
rect 1613 432 1615 452
rect 725 413 739 415
rect 725 405 739 407
rect 188 375 190 395
rect 287 389 307 391
rect 725 397 739 399
rect 725 389 739 391
rect 287 381 307 383
rect 715 317 735 319
rect 715 309 735 311
rect 715 301 735 303
rect 715 293 735 295
rect 715 285 735 287
rect 715 277 735 279
rect 1480 142 1482 162
rect 1488 142 1490 162
rect 1510 142 1512 162
rect 1518 142 1520 162
rect 1550 145 1552 165
rect 1573 158 1575 178
rect 1613 142 1615 162
rect 55 46 57 66
rect 63 46 65 66
rect 85 46 87 66
rect 93 46 95 66
rect 125 49 127 69
rect 148 62 150 82
rect 188 46 190 66
<< ndiffusion >>
rect 58 2081 59 2091
rect 61 2081 62 2091
rect 88 2081 89 2091
rect 91 2081 92 2091
rect 96 2081 97 2091
rect 99 2081 100 2091
rect 151 2077 152 2087
rect 154 2077 155 2087
rect 159 2077 160 2087
rect 162 2077 163 2087
rect 191 2080 192 2090
rect 194 2080 195 2090
rect 306 2098 307 2108
rect 309 2098 310 2108
rect 329 2092 330 2102
rect 332 2092 333 2102
rect 751 2102 771 2103
rect 751 2099 771 2100
rect 751 2094 771 2095
rect 751 2091 771 2092
rect 282 2060 283 2070
rect 285 2060 286 2070
rect 1190 2080 1191 2090
rect 1193 2080 1194 2090
rect 1213 2074 1214 2084
rect 1216 2074 1217 2084
rect 1166 2042 1167 2052
rect 1169 2042 1170 2052
rect 1479 2032 1480 2042
rect 1482 2032 1483 2042
rect 1509 2032 1510 2042
rect 1512 2032 1513 2042
rect 1517 2032 1518 2042
rect 1520 2032 1521 2042
rect 1572 2028 1573 2038
rect 1575 2028 1576 2038
rect 1580 2028 1581 2038
rect 1583 2028 1584 2038
rect 1612 2031 1613 2041
rect 1615 2031 1616 2041
rect 847 2005 867 2006
rect 847 2002 867 2003
rect 847 1997 867 1998
rect 847 1994 867 1995
rect 323 1982 343 1983
rect 323 1979 343 1980
rect 323 1974 343 1975
rect 323 1971 343 1972
rect 56 1943 57 1953
rect 59 1943 60 1953
rect 86 1943 87 1953
rect 89 1943 90 1953
rect 94 1943 95 1953
rect 97 1943 98 1953
rect 384 1961 385 1971
rect 387 1961 388 1971
rect 149 1939 150 1949
rect 152 1939 153 1949
rect 157 1939 158 1949
rect 160 1939 161 1949
rect 189 1942 190 1952
rect 192 1942 193 1952
rect 748 1841 768 1842
rect 748 1838 768 1839
rect 748 1833 768 1834
rect 748 1830 768 1831
rect 56 1802 57 1812
rect 59 1802 60 1812
rect 86 1802 87 1812
rect 89 1802 90 1812
rect 94 1802 95 1812
rect 97 1802 98 1812
rect 149 1798 150 1808
rect 152 1798 153 1808
rect 157 1798 158 1808
rect 160 1798 161 1808
rect 189 1801 190 1811
rect 192 1801 193 1811
rect 306 1815 307 1825
rect 309 1815 310 1825
rect 329 1809 330 1819
rect 332 1809 333 1819
rect 934 1820 964 1821
rect 934 1817 964 1818
rect 934 1812 964 1813
rect 934 1809 964 1810
rect 934 1804 964 1805
rect 934 1801 964 1802
rect 282 1777 283 1787
rect 285 1777 286 1787
rect 742 1775 772 1776
rect 742 1772 772 1773
rect 1188 1784 1189 1794
rect 1191 1784 1192 1794
rect 1211 1778 1212 1788
rect 1214 1778 1215 1788
rect 1479 1770 1480 1780
rect 1482 1770 1483 1780
rect 1509 1770 1510 1780
rect 1512 1770 1513 1780
rect 1517 1770 1518 1780
rect 1520 1770 1521 1780
rect 742 1767 772 1768
rect 742 1764 772 1765
rect 742 1759 772 1760
rect 742 1756 772 1757
rect 1572 1766 1573 1776
rect 1575 1766 1576 1776
rect 1580 1766 1581 1776
rect 1583 1766 1584 1776
rect 1612 1769 1613 1779
rect 1615 1769 1616 1779
rect 1164 1746 1165 1756
rect 1167 1746 1168 1756
rect 323 1699 343 1700
rect 323 1696 343 1697
rect 323 1691 343 1692
rect 323 1688 343 1689
rect 56 1660 57 1670
rect 59 1660 60 1670
rect 86 1660 87 1670
rect 89 1660 90 1670
rect 94 1660 95 1670
rect 97 1660 98 1670
rect 387 1673 388 1683
rect 390 1673 391 1683
rect 149 1656 150 1666
rect 152 1656 153 1666
rect 157 1656 158 1666
rect 160 1656 161 1666
rect 189 1659 190 1669
rect 192 1659 193 1669
rect 756 1567 776 1568
rect 756 1564 776 1565
rect 756 1559 776 1560
rect 756 1556 776 1557
rect 750 1501 780 1502
rect 56 1473 57 1483
rect 59 1473 60 1483
rect 86 1473 87 1483
rect 89 1473 90 1483
rect 94 1473 95 1483
rect 97 1473 98 1483
rect 149 1469 150 1479
rect 152 1469 153 1479
rect 157 1469 158 1479
rect 160 1469 161 1479
rect 189 1472 190 1482
rect 192 1472 193 1482
rect 306 1486 307 1496
rect 309 1486 310 1496
rect 750 1498 780 1499
rect 750 1493 780 1494
rect 329 1480 330 1490
rect 332 1480 333 1490
rect 750 1490 780 1491
rect 943 1489 983 1490
rect 750 1485 780 1486
rect 750 1482 780 1483
rect 943 1486 983 1487
rect 943 1481 983 1482
rect 943 1478 983 1479
rect 943 1473 983 1474
rect 943 1470 983 1471
rect 943 1465 983 1466
rect 943 1462 983 1463
rect 282 1448 283 1458
rect 285 1448 286 1458
rect 750 1419 790 1420
rect 750 1416 790 1417
rect 750 1411 790 1412
rect 1188 1424 1189 1434
rect 1191 1424 1192 1434
rect 1211 1418 1212 1428
rect 1214 1418 1215 1428
rect 750 1408 790 1409
rect 750 1403 790 1404
rect 750 1400 790 1401
rect 1479 1403 1480 1413
rect 1482 1403 1483 1413
rect 1509 1403 1510 1413
rect 1512 1403 1513 1413
rect 1517 1403 1518 1413
rect 1520 1403 1521 1413
rect 1572 1399 1573 1409
rect 1575 1399 1576 1409
rect 1580 1399 1581 1409
rect 1583 1399 1584 1409
rect 1612 1402 1613 1412
rect 1615 1402 1616 1412
rect 750 1395 790 1396
rect 750 1392 790 1393
rect 1164 1386 1165 1396
rect 1167 1386 1168 1396
rect 323 1370 343 1371
rect 323 1367 343 1368
rect 323 1362 343 1363
rect 323 1359 343 1360
rect 56 1331 57 1341
rect 59 1331 60 1341
rect 86 1331 87 1341
rect 89 1331 90 1341
rect 94 1331 95 1341
rect 97 1331 98 1341
rect 387 1347 388 1357
rect 390 1347 391 1357
rect 149 1327 150 1337
rect 152 1327 153 1337
rect 157 1327 158 1337
rect 160 1327 161 1337
rect 189 1330 190 1340
rect 192 1330 193 1340
rect 758 1153 778 1154
rect 758 1150 778 1151
rect 758 1145 778 1146
rect 758 1142 778 1143
rect 752 1087 782 1088
rect 752 1084 782 1085
rect 752 1079 782 1080
rect 752 1076 782 1077
rect 752 1071 782 1072
rect 752 1068 782 1069
rect 968 1034 1018 1035
rect 968 1031 1018 1032
rect 968 1026 1018 1027
rect 968 1023 1018 1024
rect 968 1018 1018 1019
rect 56 983 57 993
rect 59 983 60 993
rect 86 983 87 993
rect 89 983 90 993
rect 94 983 95 993
rect 97 983 98 993
rect 149 979 150 989
rect 152 979 153 989
rect 157 979 158 989
rect 160 979 161 989
rect 189 982 190 992
rect 192 982 193 992
rect 304 997 305 1007
rect 307 997 308 1007
rect 968 1015 1018 1016
rect 968 1010 1018 1011
rect 752 1005 792 1006
rect 327 991 328 1001
rect 330 991 331 1001
rect 752 1002 792 1003
rect 968 1007 1018 1008
rect 968 1002 1018 1003
rect 752 997 792 998
rect 968 999 1018 1000
rect 1188 1009 1189 1019
rect 1191 1009 1192 1019
rect 1211 1003 1212 1013
rect 1214 1003 1215 1013
rect 752 994 792 995
rect 752 989 792 990
rect 752 986 792 987
rect 752 981 792 982
rect 1479 985 1480 995
rect 1482 985 1483 995
rect 1509 985 1510 995
rect 1512 985 1513 995
rect 1517 985 1518 995
rect 1520 985 1521 995
rect 1572 981 1573 991
rect 1575 981 1576 991
rect 1580 981 1581 991
rect 1583 981 1584 991
rect 1612 984 1613 994
rect 1615 984 1616 994
rect 752 978 792 979
rect 1164 971 1165 981
rect 1167 971 1168 981
rect 280 959 281 969
rect 283 959 284 969
rect 753 918 803 919
rect 753 915 803 916
rect 753 910 803 911
rect 753 907 803 908
rect 753 902 803 903
rect 753 899 803 900
rect 753 894 803 895
rect 753 891 803 892
rect 753 886 803 887
rect 321 881 341 882
rect 321 878 341 879
rect 321 873 341 874
rect 753 883 803 884
rect 321 870 341 871
rect 54 842 55 852
rect 57 842 58 852
rect 84 842 85 852
rect 87 842 88 852
rect 92 842 93 852
rect 95 842 96 852
rect 386 862 387 872
rect 389 862 390 872
rect 147 838 148 848
rect 150 838 151 848
rect 155 838 156 848
rect 158 838 159 848
rect 187 841 188 851
rect 190 841 191 851
rect 757 658 777 659
rect 757 655 777 656
rect 757 650 777 651
rect 757 647 777 648
rect 751 592 781 593
rect 751 589 781 590
rect 751 584 781 585
rect 751 581 781 582
rect 751 576 781 577
rect 751 573 781 574
rect 975 526 1035 527
rect 54 493 55 503
rect 57 493 58 503
rect 84 493 85 503
rect 87 493 88 503
rect 92 493 93 503
rect 95 493 96 503
rect 147 489 148 499
rect 150 489 151 499
rect 155 489 156 499
rect 158 489 159 499
rect 187 492 188 502
rect 190 492 191 502
rect 303 507 304 517
rect 306 507 307 517
rect 975 523 1035 524
rect 975 518 1035 519
rect 326 501 327 511
rect 329 501 330 511
rect 751 510 791 511
rect 975 515 1035 516
rect 975 510 1035 511
rect 751 507 791 508
rect 751 502 791 503
rect 975 507 1035 508
rect 975 502 1035 503
rect 751 499 791 500
rect 751 494 791 495
rect 975 499 1035 500
rect 975 494 1035 495
rect 751 491 791 492
rect 751 486 791 487
rect 975 491 1035 492
rect 975 486 1035 487
rect 751 483 791 484
rect 975 483 1035 484
rect 279 469 280 479
rect 282 469 283 479
rect 1188 469 1189 479
rect 1191 469 1192 479
rect 1211 463 1212 473
rect 1214 463 1215 473
rect 1164 431 1165 441
rect 1167 431 1168 441
rect 752 423 802 424
rect 752 420 802 421
rect 752 415 802 416
rect 752 412 802 413
rect 1479 409 1480 419
rect 1482 409 1483 419
rect 1509 409 1510 419
rect 1512 409 1513 419
rect 1517 409 1518 419
rect 1520 409 1521 419
rect 752 407 802 408
rect 1572 405 1573 415
rect 1575 405 1576 415
rect 1580 405 1581 415
rect 1583 405 1584 415
rect 1612 408 1613 418
rect 1615 408 1616 418
rect 320 391 340 392
rect 320 388 340 389
rect 752 404 802 405
rect 752 399 802 400
rect 752 396 802 397
rect 752 391 802 392
rect 320 383 340 384
rect 320 380 340 381
rect 386 376 387 386
rect 389 376 390 386
rect 752 388 802 389
rect 54 352 55 362
rect 57 352 58 362
rect 84 352 85 362
rect 87 352 88 362
rect 92 352 93 362
rect 95 352 96 362
rect 147 348 148 358
rect 150 348 151 358
rect 155 348 156 358
rect 158 348 159 358
rect 187 351 188 361
rect 190 351 191 361
rect 748 319 808 320
rect 748 316 808 317
rect 748 311 808 312
rect 748 308 808 309
rect 748 303 808 304
rect 748 300 808 301
rect 748 295 808 296
rect 748 292 808 293
rect 748 287 808 288
rect 748 284 808 285
rect 748 279 808 280
rect 748 276 808 277
rect 1479 119 1480 129
rect 1482 119 1483 129
rect 1509 119 1510 129
rect 1512 119 1513 129
rect 1517 119 1518 129
rect 1520 119 1521 129
rect 1572 115 1573 125
rect 1575 115 1576 125
rect 1580 115 1581 125
rect 1583 115 1584 125
rect 1612 118 1613 128
rect 1615 118 1616 128
rect 54 23 55 33
rect 57 23 58 33
rect 84 23 85 33
rect 87 23 88 33
rect 92 23 93 33
rect 95 23 96 33
rect 147 19 148 29
rect 150 19 151 29
rect 155 19 156 29
rect 158 19 159 29
rect 187 22 188 32
rect 190 22 191 32
<< pdiffusion >>
rect 58 2104 59 2124
rect 61 2104 62 2124
rect 66 2104 67 2124
rect 69 2104 70 2124
rect 88 2104 89 2124
rect 91 2104 92 2124
rect 96 2104 97 2124
rect 99 2104 100 2124
rect 128 2107 129 2127
rect 131 2107 132 2127
rect 151 2120 152 2140
rect 154 2120 155 2140
rect 191 2104 192 2124
rect 194 2104 195 2124
rect 306 2121 307 2141
rect 309 2121 310 2141
rect 329 2121 330 2141
rect 332 2121 333 2141
rect 282 2084 283 2104
rect 285 2084 286 2104
rect 718 2102 738 2103
rect 1190 2103 1191 2123
rect 1193 2103 1194 2123
rect 1213 2103 1214 2123
rect 1216 2103 1217 2123
rect 718 2099 738 2100
rect 718 2094 738 2095
rect 718 2091 738 2092
rect 1166 2066 1167 2086
rect 1169 2066 1170 2086
rect 1479 2055 1480 2075
rect 1482 2055 1483 2075
rect 1487 2055 1488 2075
rect 1490 2055 1491 2075
rect 1509 2055 1510 2075
rect 1512 2055 1513 2075
rect 1517 2055 1518 2075
rect 1520 2055 1521 2075
rect 1549 2058 1550 2078
rect 1552 2058 1553 2078
rect 1572 2071 1573 2091
rect 1575 2071 1576 2091
rect 1612 2055 1613 2075
rect 1615 2055 1616 2075
rect 56 1966 57 1986
rect 59 1966 60 1986
rect 64 1966 65 1986
rect 67 1966 68 1986
rect 86 1966 87 1986
rect 89 1966 90 1986
rect 94 1966 95 1986
rect 97 1966 98 1986
rect 126 1969 127 1989
rect 129 1969 130 1989
rect 149 1982 150 2002
rect 152 1982 153 2002
rect 189 1966 190 1986
rect 192 1966 193 1986
rect 290 1982 310 1983
rect 384 1985 385 2005
rect 387 1985 388 2005
rect 814 2005 834 2006
rect 814 2002 834 2003
rect 814 1997 834 1998
rect 814 1994 834 1995
rect 290 1979 310 1980
rect 290 1974 310 1975
rect 290 1971 310 1972
rect 56 1825 57 1845
rect 59 1825 60 1845
rect 64 1825 65 1845
rect 67 1825 68 1845
rect 86 1825 87 1845
rect 89 1825 90 1845
rect 94 1825 95 1845
rect 97 1825 98 1845
rect 126 1828 127 1848
rect 129 1828 130 1848
rect 149 1841 150 1861
rect 152 1841 153 1861
rect 189 1825 190 1845
rect 192 1825 193 1845
rect 306 1838 307 1858
rect 309 1838 310 1858
rect 329 1838 330 1858
rect 332 1838 333 1858
rect 715 1841 735 1842
rect 715 1838 735 1839
rect 715 1833 735 1834
rect 715 1830 735 1831
rect 282 1801 283 1821
rect 285 1801 286 1821
rect 901 1820 921 1821
rect 901 1817 921 1818
rect 901 1812 921 1813
rect 901 1809 921 1810
rect 901 1804 921 1805
rect 1188 1807 1189 1827
rect 1191 1807 1192 1827
rect 1211 1807 1212 1827
rect 1214 1807 1215 1827
rect 901 1801 921 1802
rect 709 1775 729 1776
rect 709 1772 729 1773
rect 709 1767 729 1768
rect 1164 1770 1165 1790
rect 1167 1770 1168 1790
rect 1479 1793 1480 1813
rect 1482 1793 1483 1813
rect 1487 1793 1488 1813
rect 1490 1793 1491 1813
rect 1509 1793 1510 1813
rect 1512 1793 1513 1813
rect 1517 1793 1518 1813
rect 1520 1793 1521 1813
rect 1549 1796 1550 1816
rect 1552 1796 1553 1816
rect 1572 1809 1573 1829
rect 1575 1809 1576 1829
rect 1612 1793 1613 1813
rect 1615 1793 1616 1813
rect 709 1764 729 1765
rect 709 1759 729 1760
rect 709 1756 729 1757
rect 56 1683 57 1703
rect 59 1683 60 1703
rect 64 1683 65 1703
rect 67 1683 68 1703
rect 86 1683 87 1703
rect 89 1683 90 1703
rect 94 1683 95 1703
rect 97 1683 98 1703
rect 126 1686 127 1706
rect 129 1686 130 1706
rect 149 1699 150 1719
rect 152 1699 153 1719
rect 189 1683 190 1703
rect 192 1683 193 1703
rect 290 1699 310 1700
rect 387 1697 388 1717
rect 390 1697 391 1717
rect 290 1696 310 1697
rect 290 1691 310 1692
rect 290 1688 310 1689
rect 723 1567 743 1568
rect 723 1564 743 1565
rect 723 1559 743 1560
rect 723 1556 743 1557
rect 56 1496 57 1516
rect 59 1496 60 1516
rect 64 1496 65 1516
rect 67 1496 68 1516
rect 86 1496 87 1516
rect 89 1496 90 1516
rect 94 1496 95 1516
rect 97 1496 98 1516
rect 126 1499 127 1519
rect 129 1499 130 1519
rect 149 1512 150 1532
rect 152 1512 153 1532
rect 189 1496 190 1516
rect 192 1496 193 1516
rect 306 1509 307 1529
rect 309 1509 310 1529
rect 329 1509 330 1529
rect 332 1509 333 1529
rect 717 1501 737 1502
rect 717 1498 737 1499
rect 282 1472 283 1492
rect 285 1472 286 1492
rect 717 1493 737 1494
rect 717 1490 737 1491
rect 717 1485 737 1486
rect 910 1489 930 1490
rect 910 1486 930 1487
rect 717 1482 737 1483
rect 910 1481 930 1482
rect 910 1478 930 1479
rect 910 1473 930 1474
rect 910 1470 930 1471
rect 910 1465 930 1466
rect 910 1462 930 1463
rect 1188 1447 1189 1467
rect 1191 1447 1192 1467
rect 1211 1447 1212 1467
rect 1214 1447 1215 1467
rect 717 1419 737 1420
rect 717 1416 737 1417
rect 717 1411 737 1412
rect 1164 1410 1165 1430
rect 1167 1410 1168 1430
rect 1479 1426 1480 1446
rect 1482 1426 1483 1446
rect 1487 1426 1488 1446
rect 1490 1426 1491 1446
rect 1509 1426 1510 1446
rect 1512 1426 1513 1446
rect 1517 1426 1518 1446
rect 1520 1426 1521 1446
rect 1549 1429 1550 1449
rect 1552 1429 1553 1449
rect 1572 1442 1573 1462
rect 1575 1442 1576 1462
rect 1612 1426 1613 1446
rect 1615 1426 1616 1446
rect 717 1408 737 1409
rect 717 1403 737 1404
rect 717 1400 737 1401
rect 717 1395 737 1396
rect 717 1392 737 1393
rect 56 1354 57 1374
rect 59 1354 60 1374
rect 64 1354 65 1374
rect 67 1354 68 1374
rect 86 1354 87 1374
rect 89 1354 90 1374
rect 94 1354 95 1374
rect 97 1354 98 1374
rect 126 1357 127 1377
rect 129 1357 130 1377
rect 149 1370 150 1390
rect 152 1370 153 1390
rect 189 1354 190 1374
rect 192 1354 193 1374
rect 290 1370 310 1371
rect 387 1371 388 1391
rect 390 1371 391 1391
rect 290 1367 310 1368
rect 290 1362 310 1363
rect 290 1359 310 1360
rect 725 1153 745 1154
rect 725 1150 745 1151
rect 725 1145 745 1146
rect 725 1142 745 1143
rect 719 1087 739 1088
rect 719 1084 739 1085
rect 719 1079 739 1080
rect 719 1076 739 1077
rect 719 1071 739 1072
rect 719 1068 739 1069
rect 56 1006 57 1026
rect 59 1006 60 1026
rect 64 1006 65 1026
rect 67 1006 68 1026
rect 86 1006 87 1026
rect 89 1006 90 1026
rect 94 1006 95 1026
rect 97 1006 98 1026
rect 126 1009 127 1029
rect 129 1009 130 1029
rect 149 1022 150 1042
rect 152 1022 153 1042
rect 189 1006 190 1026
rect 192 1006 193 1026
rect 304 1020 305 1040
rect 307 1020 308 1040
rect 327 1020 328 1040
rect 330 1020 331 1040
rect 941 1034 955 1035
rect 1188 1032 1189 1052
rect 1191 1032 1192 1052
rect 1211 1032 1212 1052
rect 1214 1032 1215 1052
rect 941 1031 955 1032
rect 941 1026 955 1027
rect 941 1023 955 1024
rect 941 1018 955 1019
rect 941 1015 955 1016
rect 280 983 281 1003
rect 283 983 284 1003
rect 719 1005 739 1006
rect 941 1010 955 1011
rect 941 1007 955 1008
rect 719 1002 739 1003
rect 719 997 739 998
rect 941 1002 955 1003
rect 941 999 955 1000
rect 1164 995 1165 1015
rect 1167 995 1168 1015
rect 1479 1008 1480 1028
rect 1482 1008 1483 1028
rect 1487 1008 1488 1028
rect 1490 1008 1491 1028
rect 1509 1008 1510 1028
rect 1512 1008 1513 1028
rect 1517 1008 1518 1028
rect 1520 1008 1521 1028
rect 1549 1011 1550 1031
rect 1552 1011 1553 1031
rect 1572 1024 1573 1044
rect 1575 1024 1576 1044
rect 1612 1008 1613 1028
rect 1615 1008 1616 1028
rect 719 994 739 995
rect 719 989 739 990
rect 719 986 739 987
rect 719 981 739 982
rect 719 978 739 979
rect 726 918 740 919
rect 726 915 740 916
rect 726 910 740 911
rect 726 907 740 908
rect 54 865 55 885
rect 57 865 58 885
rect 62 865 63 885
rect 65 865 66 885
rect 84 865 85 885
rect 87 865 88 885
rect 92 865 93 885
rect 95 865 96 885
rect 124 868 125 888
rect 127 868 128 888
rect 147 881 148 901
rect 150 881 151 901
rect 386 886 387 906
rect 389 886 390 906
rect 726 902 740 903
rect 726 899 740 900
rect 726 894 740 895
rect 726 891 740 892
rect 726 886 740 887
rect 187 865 188 885
rect 190 865 191 885
rect 288 881 308 882
rect 288 878 308 879
rect 288 873 308 874
rect 726 883 740 884
rect 288 870 308 871
rect 724 658 744 659
rect 724 655 744 656
rect 724 650 744 651
rect 724 647 744 648
rect 718 592 738 593
rect 718 589 738 590
rect 718 584 738 585
rect 718 581 738 582
rect 718 576 738 577
rect 718 573 738 574
rect 54 516 55 536
rect 57 516 58 536
rect 62 516 63 536
rect 65 516 66 536
rect 84 516 85 536
rect 87 516 88 536
rect 92 516 93 536
rect 95 516 96 536
rect 124 519 125 539
rect 127 519 128 539
rect 147 532 148 552
rect 150 532 151 552
rect 187 516 188 536
rect 190 516 191 536
rect 303 530 304 550
rect 306 530 307 550
rect 326 530 327 550
rect 329 530 330 550
rect 942 526 962 527
rect 942 523 962 524
rect 279 493 280 513
rect 282 493 283 513
rect 942 518 962 519
rect 942 515 962 516
rect 718 510 738 511
rect 942 510 962 511
rect 718 507 738 508
rect 718 502 738 503
rect 942 507 962 508
rect 942 502 962 503
rect 718 499 738 500
rect 718 494 738 495
rect 942 499 962 500
rect 942 494 962 495
rect 1188 492 1189 512
rect 1191 492 1192 512
rect 1211 492 1212 512
rect 1214 492 1215 512
rect 718 491 738 492
rect 718 486 738 487
rect 942 491 962 492
rect 942 486 962 487
rect 718 483 738 484
rect 942 483 962 484
rect 1164 455 1165 475
rect 1167 455 1168 475
rect 1479 432 1480 452
rect 1482 432 1483 452
rect 1487 432 1488 452
rect 1490 432 1491 452
rect 1509 432 1510 452
rect 1512 432 1513 452
rect 1517 432 1518 452
rect 1520 432 1521 452
rect 1549 435 1550 455
rect 1552 435 1553 455
rect 1572 448 1573 468
rect 1575 448 1576 468
rect 725 423 739 424
rect 725 420 739 421
rect 54 375 55 395
rect 57 375 58 395
rect 62 375 63 395
rect 65 375 66 395
rect 84 375 85 395
rect 87 375 88 395
rect 92 375 93 395
rect 95 375 96 395
rect 124 378 125 398
rect 127 378 128 398
rect 147 391 148 411
rect 150 391 151 411
rect 386 400 387 420
rect 389 400 390 420
rect 725 415 739 416
rect 1612 432 1613 452
rect 1615 432 1616 452
rect 725 412 739 413
rect 725 407 739 408
rect 725 404 739 405
rect 187 375 188 395
rect 190 375 191 395
rect 287 391 307 392
rect 287 388 307 389
rect 287 383 307 384
rect 725 399 739 400
rect 725 396 739 397
rect 725 391 739 392
rect 725 388 739 389
rect 287 380 307 381
rect 715 319 735 320
rect 715 316 735 317
rect 715 311 735 312
rect 715 308 735 309
rect 715 303 735 304
rect 715 300 735 301
rect 715 295 735 296
rect 715 292 735 293
rect 715 287 735 288
rect 715 284 735 285
rect 715 279 735 280
rect 715 276 735 277
rect 1479 142 1480 162
rect 1482 142 1483 162
rect 1487 142 1488 162
rect 1490 142 1491 162
rect 1509 142 1510 162
rect 1512 142 1513 162
rect 1517 142 1518 162
rect 1520 142 1521 162
rect 1549 145 1550 165
rect 1552 145 1553 165
rect 1572 158 1573 178
rect 1575 158 1576 178
rect 1612 142 1613 162
rect 1615 142 1616 162
rect 54 46 55 66
rect 57 46 58 66
rect 62 46 63 66
rect 65 46 66 66
rect 84 46 85 66
rect 87 46 88 66
rect 92 46 93 66
rect 95 46 96 66
rect 124 49 125 69
rect 127 49 128 69
rect 147 62 148 82
rect 150 62 151 82
rect 187 46 188 66
rect 190 46 191 66
<< ndcontact >>
rect 54 2081 58 2091
rect 62 2081 74 2091
rect 84 2081 88 2091
rect 92 2081 96 2091
rect 100 2081 104 2091
rect 147 2077 151 2087
rect 155 2077 159 2087
rect 163 2077 167 2087
rect 187 2080 191 2090
rect 195 2080 199 2090
rect 302 2098 306 2108
rect 310 2098 314 2108
rect 325 2092 329 2102
rect 333 2092 337 2102
rect 751 2103 771 2107
rect 751 2095 771 2099
rect 751 2087 771 2091
rect 278 2060 282 2070
rect 286 2060 290 2070
rect 1186 2080 1190 2090
rect 1194 2080 1198 2090
rect 1209 2074 1213 2084
rect 1217 2074 1221 2084
rect 1162 2042 1166 2052
rect 1170 2042 1174 2052
rect 1475 2032 1479 2042
rect 1483 2032 1495 2042
rect 1505 2032 1509 2042
rect 1513 2032 1517 2042
rect 1521 2032 1525 2042
rect 1568 2028 1572 2038
rect 1576 2028 1580 2038
rect 1584 2028 1588 2038
rect 1608 2031 1612 2041
rect 1616 2031 1620 2041
rect 323 1983 343 1987
rect 847 2006 867 2010
rect 847 1998 867 2002
rect 847 1990 867 1994
rect 323 1975 343 1979
rect 323 1967 343 1971
rect 52 1943 56 1953
rect 60 1943 72 1953
rect 82 1943 86 1953
rect 90 1943 94 1953
rect 98 1943 102 1953
rect 380 1961 384 1971
rect 388 1961 392 1971
rect 145 1939 149 1949
rect 153 1939 157 1949
rect 161 1939 165 1949
rect 185 1942 189 1952
rect 193 1942 197 1952
rect 748 1842 768 1846
rect 748 1834 768 1838
rect 748 1826 768 1830
rect 52 1802 56 1812
rect 60 1802 72 1812
rect 82 1802 86 1812
rect 90 1802 94 1812
rect 98 1802 102 1812
rect 145 1798 149 1808
rect 153 1798 157 1808
rect 161 1798 165 1808
rect 185 1801 189 1811
rect 193 1801 197 1811
rect 302 1815 306 1825
rect 310 1815 314 1825
rect 325 1809 329 1819
rect 333 1809 337 1819
rect 934 1821 964 1825
rect 934 1813 964 1817
rect 934 1805 964 1809
rect 934 1797 964 1801
rect 278 1777 282 1787
rect 286 1777 290 1787
rect 742 1776 772 1780
rect 742 1768 772 1772
rect 1184 1784 1188 1794
rect 1192 1784 1196 1794
rect 1207 1778 1211 1788
rect 1215 1778 1219 1788
rect 1475 1770 1479 1780
rect 1483 1770 1495 1780
rect 1505 1770 1509 1780
rect 1513 1770 1517 1780
rect 1521 1770 1525 1780
rect 742 1760 772 1764
rect 1568 1766 1572 1776
rect 1576 1766 1580 1776
rect 1584 1766 1588 1776
rect 1608 1769 1612 1779
rect 1616 1769 1620 1779
rect 742 1752 772 1756
rect 1160 1746 1164 1756
rect 1168 1746 1172 1756
rect 323 1700 343 1704
rect 323 1692 343 1696
rect 323 1684 343 1688
rect 52 1660 56 1670
rect 60 1660 72 1670
rect 82 1660 86 1670
rect 90 1660 94 1670
rect 98 1660 102 1670
rect 383 1673 387 1683
rect 391 1673 395 1683
rect 145 1656 149 1666
rect 153 1656 157 1666
rect 161 1656 165 1666
rect 185 1659 189 1669
rect 193 1659 197 1669
rect 756 1568 776 1572
rect 756 1560 776 1564
rect 756 1552 776 1556
rect 750 1502 780 1506
rect 52 1473 56 1483
rect 60 1473 72 1483
rect 82 1473 86 1483
rect 90 1473 94 1483
rect 98 1473 102 1483
rect 145 1469 149 1479
rect 153 1469 157 1479
rect 161 1469 165 1479
rect 185 1472 189 1482
rect 193 1472 197 1482
rect 302 1486 306 1496
rect 310 1486 314 1496
rect 750 1494 780 1498
rect 325 1480 329 1490
rect 333 1480 337 1490
rect 750 1486 780 1490
rect 943 1490 983 1494
rect 750 1478 780 1482
rect 943 1482 983 1486
rect 943 1474 983 1478
rect 943 1466 983 1470
rect 943 1458 983 1462
rect 278 1448 282 1458
rect 286 1448 290 1458
rect 750 1420 790 1424
rect 750 1412 790 1416
rect 1184 1424 1188 1434
rect 1192 1424 1196 1434
rect 1207 1418 1211 1428
rect 1215 1418 1219 1428
rect 750 1404 790 1408
rect 750 1396 790 1400
rect 1475 1403 1479 1413
rect 1483 1403 1495 1413
rect 1505 1403 1509 1413
rect 1513 1403 1517 1413
rect 1521 1403 1525 1413
rect 1568 1399 1572 1409
rect 1576 1399 1580 1409
rect 1584 1399 1588 1409
rect 1608 1402 1612 1412
rect 1616 1402 1620 1412
rect 323 1371 343 1375
rect 750 1388 790 1392
rect 1160 1386 1164 1396
rect 1168 1386 1172 1396
rect 323 1363 343 1367
rect 323 1355 343 1359
rect 52 1331 56 1341
rect 60 1331 72 1341
rect 82 1331 86 1341
rect 90 1331 94 1341
rect 98 1331 102 1341
rect 383 1347 387 1357
rect 391 1347 395 1357
rect 145 1327 149 1337
rect 153 1327 157 1337
rect 161 1327 165 1337
rect 185 1330 189 1340
rect 193 1330 197 1340
rect 758 1154 778 1158
rect 758 1146 778 1150
rect 758 1138 778 1142
rect 752 1088 782 1092
rect 752 1080 782 1084
rect 752 1072 782 1076
rect 752 1064 782 1068
rect 968 1035 1018 1039
rect 968 1027 1018 1031
rect 968 1019 1018 1023
rect 52 983 56 993
rect 60 983 72 993
rect 82 983 86 993
rect 90 983 94 993
rect 98 983 102 993
rect 145 979 149 989
rect 153 979 157 989
rect 161 979 165 989
rect 185 982 189 992
rect 193 982 197 992
rect 300 997 304 1007
rect 308 997 312 1007
rect 752 1006 792 1010
rect 968 1011 1018 1015
rect 323 991 327 1001
rect 331 991 335 1001
rect 752 998 792 1002
rect 968 1003 1018 1007
rect 968 995 1018 999
rect 1184 1009 1188 1019
rect 1192 1009 1196 1019
rect 1207 1003 1211 1013
rect 1215 1003 1219 1013
rect 752 990 792 994
rect 752 982 792 986
rect 1475 985 1479 995
rect 1483 985 1495 995
rect 1505 985 1509 995
rect 1513 985 1517 995
rect 1521 985 1525 995
rect 1568 981 1572 991
rect 1576 981 1580 991
rect 1584 981 1588 991
rect 1608 984 1612 994
rect 1616 984 1620 994
rect 752 974 792 978
rect 1160 971 1164 981
rect 1168 971 1172 981
rect 276 959 280 969
rect 284 959 288 969
rect 753 919 803 923
rect 753 911 803 915
rect 753 903 803 907
rect 753 895 803 899
rect 753 887 803 891
rect 321 882 341 886
rect 321 874 341 878
rect 753 879 803 883
rect 321 866 341 870
rect 50 842 54 852
rect 58 842 70 852
rect 80 842 84 852
rect 88 842 92 852
rect 96 842 100 852
rect 382 862 386 872
rect 390 862 394 872
rect 143 838 147 848
rect 151 838 155 848
rect 159 838 163 848
rect 183 841 187 851
rect 191 841 195 851
rect 757 659 777 663
rect 757 651 777 655
rect 757 643 777 647
rect 751 593 781 597
rect 751 585 781 589
rect 751 577 781 581
rect 751 569 781 573
rect 975 527 1035 531
rect 50 493 54 503
rect 58 493 70 503
rect 80 493 84 503
rect 88 493 92 503
rect 96 493 100 503
rect 143 489 147 499
rect 151 489 155 499
rect 159 489 163 499
rect 183 492 187 502
rect 191 492 195 502
rect 299 507 303 517
rect 307 507 311 517
rect 975 519 1035 523
rect 322 501 326 511
rect 330 501 334 511
rect 751 511 791 515
rect 975 511 1035 515
rect 751 503 791 507
rect 975 503 1035 507
rect 751 495 791 499
rect 975 495 1035 499
rect 751 487 791 491
rect 975 487 1035 491
rect 751 479 791 483
rect 975 479 1035 483
rect 275 469 279 479
rect 283 469 287 479
rect 1184 469 1188 479
rect 1192 469 1196 479
rect 1207 463 1211 473
rect 1215 463 1219 473
rect 1160 431 1164 441
rect 1168 431 1172 441
rect 752 424 802 428
rect 752 416 802 420
rect 752 408 802 412
rect 1475 409 1479 419
rect 1483 409 1495 419
rect 1505 409 1509 419
rect 1513 409 1517 419
rect 1521 409 1525 419
rect 1568 405 1572 415
rect 1576 405 1580 415
rect 1584 405 1588 415
rect 1608 408 1612 418
rect 1616 408 1620 418
rect 320 392 340 396
rect 320 384 340 388
rect 752 400 802 404
rect 752 392 802 396
rect 320 376 340 380
rect 382 376 386 386
rect 390 376 394 386
rect 752 384 802 388
rect 50 352 54 362
rect 58 352 70 362
rect 80 352 84 362
rect 88 352 92 362
rect 96 352 100 362
rect 143 348 147 358
rect 151 348 155 358
rect 159 348 163 358
rect 183 351 187 361
rect 191 351 195 361
rect 748 320 808 324
rect 748 312 808 316
rect 748 304 808 308
rect 748 296 808 300
rect 748 288 808 292
rect 748 280 808 284
rect 748 272 808 276
rect 1475 119 1479 129
rect 1483 119 1495 129
rect 1505 119 1509 129
rect 1513 119 1517 129
rect 1521 119 1525 129
rect 1568 115 1572 125
rect 1576 115 1580 125
rect 1584 115 1588 125
rect 1608 118 1612 128
rect 1616 118 1620 128
rect 50 23 54 33
rect 58 23 70 33
rect 80 23 84 33
rect 88 23 92 33
rect 96 23 100 33
rect 143 19 147 29
rect 151 19 155 29
rect 159 19 163 29
rect 183 22 187 32
rect 191 22 195 32
<< pdcontact >>
rect 54 2104 58 2124
rect 62 2104 66 2124
rect 70 2104 74 2124
rect 84 2104 88 2124
rect 92 2104 96 2124
rect 100 2104 104 2124
rect 124 2107 128 2127
rect 132 2107 136 2127
rect 147 2120 151 2140
rect 155 2120 167 2140
rect 187 2104 191 2124
rect 195 2104 199 2124
rect 302 2121 306 2141
rect 310 2121 314 2141
rect 325 2121 329 2141
rect 333 2121 337 2141
rect 278 2084 282 2104
rect 286 2084 290 2104
rect 718 2103 738 2107
rect 1186 2103 1190 2123
rect 1194 2103 1198 2123
rect 1209 2103 1213 2123
rect 1217 2103 1221 2123
rect 718 2095 738 2099
rect 718 2087 738 2091
rect 1162 2066 1166 2086
rect 1170 2066 1174 2086
rect 1475 2055 1479 2075
rect 1483 2055 1487 2075
rect 1491 2055 1495 2075
rect 1505 2055 1509 2075
rect 1513 2055 1517 2075
rect 1521 2055 1525 2075
rect 1545 2058 1549 2078
rect 1553 2058 1557 2078
rect 1568 2071 1572 2091
rect 1576 2071 1588 2091
rect 1608 2055 1612 2075
rect 1616 2055 1620 2075
rect 52 1966 56 1986
rect 60 1966 64 1986
rect 68 1966 72 1986
rect 82 1966 86 1986
rect 90 1966 94 1986
rect 98 1966 102 1986
rect 122 1969 126 1989
rect 130 1969 134 1989
rect 145 1982 149 2002
rect 153 1982 165 2002
rect 185 1966 189 1986
rect 193 1966 197 1986
rect 290 1983 310 1987
rect 380 1985 384 2005
rect 388 1985 392 2005
rect 814 2006 834 2010
rect 814 1998 834 2002
rect 814 1990 834 1994
rect 290 1975 310 1979
rect 290 1967 310 1971
rect 52 1825 56 1845
rect 60 1825 64 1845
rect 68 1825 72 1845
rect 82 1825 86 1845
rect 90 1825 94 1845
rect 98 1825 102 1845
rect 122 1828 126 1848
rect 130 1828 134 1848
rect 145 1841 149 1861
rect 153 1841 165 1861
rect 185 1825 189 1845
rect 193 1825 197 1845
rect 302 1838 306 1858
rect 310 1838 314 1858
rect 325 1838 329 1858
rect 333 1838 337 1858
rect 715 1842 735 1846
rect 715 1834 735 1838
rect 715 1826 735 1830
rect 278 1801 282 1821
rect 286 1801 290 1821
rect 901 1821 921 1825
rect 901 1813 921 1817
rect 901 1805 921 1809
rect 1184 1807 1188 1827
rect 1192 1807 1196 1827
rect 1207 1807 1211 1827
rect 1215 1807 1219 1827
rect 901 1797 921 1801
rect 709 1776 729 1780
rect 709 1768 729 1772
rect 1160 1770 1164 1790
rect 1168 1770 1172 1790
rect 1475 1793 1479 1813
rect 1483 1793 1487 1813
rect 1491 1793 1495 1813
rect 1505 1793 1509 1813
rect 1513 1793 1517 1813
rect 1521 1793 1525 1813
rect 1545 1796 1549 1816
rect 1553 1796 1557 1816
rect 1568 1809 1572 1829
rect 1576 1809 1588 1829
rect 1608 1793 1612 1813
rect 1616 1793 1620 1813
rect 709 1760 729 1764
rect 709 1752 729 1756
rect 52 1683 56 1703
rect 60 1683 64 1703
rect 68 1683 72 1703
rect 82 1683 86 1703
rect 90 1683 94 1703
rect 98 1683 102 1703
rect 122 1686 126 1706
rect 130 1686 134 1706
rect 145 1699 149 1719
rect 153 1699 165 1719
rect 185 1683 189 1703
rect 193 1683 197 1703
rect 290 1700 310 1704
rect 383 1697 387 1717
rect 391 1697 395 1717
rect 290 1692 310 1696
rect 290 1684 310 1688
rect 723 1568 743 1572
rect 723 1560 743 1564
rect 723 1552 743 1556
rect 52 1496 56 1516
rect 60 1496 64 1516
rect 68 1496 72 1516
rect 82 1496 86 1516
rect 90 1496 94 1516
rect 98 1496 102 1516
rect 122 1499 126 1519
rect 130 1499 134 1519
rect 145 1512 149 1532
rect 153 1512 165 1532
rect 185 1496 189 1516
rect 193 1496 197 1516
rect 302 1509 306 1529
rect 310 1509 314 1529
rect 325 1509 329 1529
rect 333 1509 337 1529
rect 717 1502 737 1506
rect 278 1472 282 1492
rect 286 1472 290 1492
rect 717 1494 737 1498
rect 717 1486 737 1490
rect 910 1490 930 1494
rect 717 1478 737 1482
rect 910 1482 930 1486
rect 910 1474 930 1478
rect 910 1466 930 1470
rect 910 1458 930 1462
rect 1184 1447 1188 1467
rect 1192 1447 1196 1467
rect 1207 1447 1211 1467
rect 1215 1447 1219 1467
rect 717 1420 737 1424
rect 717 1412 737 1416
rect 1160 1410 1164 1430
rect 1168 1410 1172 1430
rect 1475 1426 1479 1446
rect 1483 1426 1487 1446
rect 1491 1426 1495 1446
rect 1505 1426 1509 1446
rect 1513 1426 1517 1446
rect 1521 1426 1525 1446
rect 1545 1429 1549 1449
rect 1553 1429 1557 1449
rect 1568 1442 1572 1462
rect 1576 1442 1588 1462
rect 1608 1426 1612 1446
rect 1616 1426 1620 1446
rect 717 1404 737 1408
rect 717 1396 737 1400
rect 52 1354 56 1374
rect 60 1354 64 1374
rect 68 1354 72 1374
rect 82 1354 86 1374
rect 90 1354 94 1374
rect 98 1354 102 1374
rect 122 1357 126 1377
rect 130 1357 134 1377
rect 145 1370 149 1390
rect 153 1370 165 1390
rect 185 1354 189 1374
rect 193 1354 197 1374
rect 290 1371 310 1375
rect 383 1371 387 1391
rect 391 1371 395 1391
rect 717 1388 737 1392
rect 290 1363 310 1367
rect 290 1355 310 1359
rect 725 1154 745 1158
rect 725 1146 745 1150
rect 725 1138 745 1142
rect 719 1088 739 1092
rect 719 1080 739 1084
rect 719 1072 739 1076
rect 719 1064 739 1068
rect 52 1006 56 1026
rect 60 1006 64 1026
rect 68 1006 72 1026
rect 82 1006 86 1026
rect 90 1006 94 1026
rect 98 1006 102 1026
rect 122 1009 126 1029
rect 130 1009 134 1029
rect 145 1022 149 1042
rect 153 1022 165 1042
rect 185 1006 189 1026
rect 193 1006 197 1026
rect 300 1020 304 1040
rect 308 1020 312 1040
rect 323 1020 327 1040
rect 331 1020 335 1040
rect 941 1035 955 1039
rect 1184 1032 1188 1052
rect 1192 1032 1196 1052
rect 1207 1032 1211 1052
rect 1215 1032 1219 1052
rect 941 1027 955 1031
rect 941 1019 955 1023
rect 941 1011 955 1015
rect 276 983 280 1003
rect 284 983 288 1003
rect 719 1006 739 1010
rect 941 1003 955 1007
rect 719 998 739 1002
rect 941 995 955 999
rect 1160 995 1164 1015
rect 1168 995 1172 1015
rect 1475 1008 1479 1028
rect 1483 1008 1487 1028
rect 1491 1008 1495 1028
rect 1505 1008 1509 1028
rect 1513 1008 1517 1028
rect 1521 1008 1525 1028
rect 1545 1011 1549 1031
rect 1553 1011 1557 1031
rect 1568 1024 1572 1044
rect 1576 1024 1588 1044
rect 1608 1008 1612 1028
rect 1616 1008 1620 1028
rect 719 990 739 994
rect 719 982 739 986
rect 719 974 739 978
rect 726 919 740 923
rect 726 911 740 915
rect 50 865 54 885
rect 58 865 62 885
rect 66 865 70 885
rect 80 865 84 885
rect 88 865 92 885
rect 96 865 100 885
rect 120 868 124 888
rect 128 868 132 888
rect 143 881 147 901
rect 151 881 163 901
rect 382 886 386 906
rect 390 886 394 906
rect 726 903 740 907
rect 726 895 740 899
rect 726 887 740 891
rect 183 865 187 885
rect 191 865 195 885
rect 288 882 308 886
rect 288 874 308 878
rect 726 879 740 883
rect 288 866 308 870
rect 724 659 744 663
rect 724 651 744 655
rect 724 643 744 647
rect 718 593 738 597
rect 718 585 738 589
rect 718 577 738 581
rect 718 569 738 573
rect 50 516 54 536
rect 58 516 62 536
rect 66 516 70 536
rect 80 516 84 536
rect 88 516 92 536
rect 96 516 100 536
rect 120 519 124 539
rect 128 519 132 539
rect 143 532 147 552
rect 151 532 163 552
rect 183 516 187 536
rect 191 516 195 536
rect 299 530 303 550
rect 307 530 311 550
rect 322 530 326 550
rect 330 530 334 550
rect 942 527 962 531
rect 275 493 279 513
rect 283 493 287 513
rect 942 519 962 523
rect 718 511 738 515
rect 942 511 962 515
rect 718 503 738 507
rect 942 503 962 507
rect 718 495 738 499
rect 942 495 962 499
rect 1184 492 1188 512
rect 1192 492 1196 512
rect 1207 492 1211 512
rect 1215 492 1219 512
rect 718 487 738 491
rect 942 487 962 491
rect 718 479 738 483
rect 942 479 962 483
rect 1160 455 1164 475
rect 1168 455 1172 475
rect 1475 432 1479 452
rect 1483 432 1487 452
rect 1491 432 1495 452
rect 1505 432 1509 452
rect 1513 432 1517 452
rect 1521 432 1525 452
rect 1545 435 1549 455
rect 1553 435 1557 455
rect 1568 448 1572 468
rect 1576 448 1588 468
rect 725 424 739 428
rect 50 375 54 395
rect 58 375 62 395
rect 66 375 70 395
rect 80 375 84 395
rect 88 375 92 395
rect 96 375 100 395
rect 120 378 124 398
rect 128 378 132 398
rect 143 391 147 411
rect 151 391 163 411
rect 382 400 386 420
rect 390 400 394 420
rect 725 416 739 420
rect 1608 432 1612 452
rect 1616 432 1620 452
rect 725 408 739 412
rect 725 400 739 404
rect 183 375 187 395
rect 191 375 195 395
rect 287 392 307 396
rect 287 384 307 388
rect 725 392 739 396
rect 287 376 307 380
rect 725 384 739 388
rect 715 320 735 324
rect 715 312 735 316
rect 715 304 735 308
rect 715 296 735 300
rect 715 288 735 292
rect 715 280 735 284
rect 715 272 735 276
rect 1475 142 1479 162
rect 1483 142 1487 162
rect 1491 142 1495 162
rect 1505 142 1509 162
rect 1513 142 1517 162
rect 1521 142 1525 162
rect 1545 145 1549 165
rect 1553 145 1557 165
rect 1568 158 1572 178
rect 1576 158 1588 178
rect 1608 142 1612 162
rect 1616 142 1620 162
rect 50 46 54 66
rect 58 46 62 66
rect 66 46 70 66
rect 80 46 84 66
rect 88 46 92 66
rect 96 46 100 66
rect 120 49 124 69
rect 128 49 132 69
rect 143 62 147 82
rect 151 62 163 82
rect 183 46 187 66
rect 191 46 195 66
<< psubstratepcontact >>
rect 42 2058 46 2063
rect 278 2052 282 2056
rect 347 1967 351 1971
rect 380 1953 384 1957
rect 40 1920 44 1925
rect 40 1779 44 1784
rect 278 1769 282 1773
rect 1160 1738 1164 1742
rect 347 1684 351 1688
rect 383 1665 387 1669
rect 40 1637 44 1642
rect 40 1450 44 1455
rect 278 1440 282 1444
rect 1160 1378 1164 1382
rect 1463 1380 1467 1385
rect 347 1355 351 1359
rect 383 1339 387 1343
rect 40 1308 44 1313
rect 40 960 44 965
rect 1160 963 1164 967
rect 1463 962 1467 967
rect 276 951 280 955
rect 345 866 349 870
rect 382 854 386 858
rect 38 819 42 824
rect 38 470 42 475
rect 275 461 279 465
rect 1160 423 1164 427
rect 344 376 348 380
rect 1463 386 1467 391
rect 382 368 386 372
rect 38 329 42 334
rect 1463 96 1467 101
rect 38 0 42 5
<< nsubstratencontact >>
rect 197 2148 201 2152
rect 278 2108 282 2112
rect 709 2087 713 2091
rect 1162 2090 1166 2094
rect 1618 2099 1622 2103
rect 195 2010 199 2014
rect 380 2009 384 2013
rect 805 1990 809 1994
rect 281 1967 285 1971
rect 195 1869 199 1873
rect 278 1825 282 1829
rect 706 1826 710 1830
rect 1618 1837 1622 1841
rect 892 1797 896 1801
rect 1160 1794 1164 1798
rect 700 1752 704 1756
rect 195 1727 199 1731
rect 383 1721 387 1725
rect 281 1684 285 1688
rect 714 1552 718 1556
rect 195 1540 199 1544
rect 278 1496 282 1500
rect 708 1478 712 1482
rect 1618 1470 1622 1474
rect 901 1458 905 1462
rect 1160 1434 1164 1438
rect 195 1398 199 1402
rect 383 1395 387 1399
rect 708 1388 712 1392
rect 281 1355 285 1359
rect 716 1138 720 1142
rect 710 1064 714 1068
rect 195 1050 199 1054
rect 1618 1052 1622 1056
rect 276 1007 280 1011
rect 1160 1019 1164 1023
rect 928 995 932 999
rect 710 974 714 978
rect 193 909 197 913
rect 382 910 386 914
rect 713 879 717 883
rect 279 866 283 870
rect 715 643 719 647
rect 709 569 713 573
rect 193 560 197 564
rect 275 517 279 521
rect 709 479 713 483
rect 933 479 937 483
rect 1160 479 1164 483
rect 1618 476 1622 480
rect 382 424 386 428
rect 193 419 197 423
rect 278 376 282 380
rect 712 384 716 388
rect 706 272 710 276
rect 1618 186 1622 190
rect 193 90 197 94
<< polysilicon >>
rect 152 2140 154 2144
rect 307 2141 309 2154
rect 330 2141 332 2145
rect 59 2124 61 2128
rect 67 2124 69 2128
rect 89 2124 91 2128
rect 97 2124 99 2128
rect 129 2127 131 2131
rect 192 2124 194 2128
rect 59 2091 61 2104
rect 67 2100 69 2104
rect 89 2091 91 2104
rect 97 2091 99 2104
rect 129 2103 131 2107
rect 152 2101 154 2120
rect 1191 2123 1193 2136
rect 1214 2123 1216 2127
rect 307 2108 309 2121
rect 330 2117 332 2121
rect 283 2104 285 2107
rect 152 2087 154 2092
rect 160 2087 162 2091
rect 192 2090 194 2104
rect 59 2077 61 2081
rect 89 2077 91 2081
rect 97 2077 99 2081
rect 330 2102 332 2109
rect 307 2095 309 2098
rect 701 2100 718 2102
rect 738 2100 751 2102
rect 771 2100 774 2102
rect 701 2092 718 2094
rect 738 2092 751 2094
rect 771 2092 774 2094
rect 330 2089 332 2092
rect 1191 2090 1193 2103
rect 1214 2099 1216 2103
rect 1573 2091 1575 2095
rect 1167 2086 1169 2089
rect 192 2077 194 2080
rect 152 2073 154 2077
rect 160 2073 162 2077
rect 283 2070 285 2084
rect 1214 2084 1216 2091
rect 1191 2077 1193 2080
rect 1480 2075 1482 2079
rect 1488 2075 1490 2079
rect 1510 2075 1512 2079
rect 1518 2075 1520 2079
rect 1550 2078 1552 2082
rect 1214 2071 1216 2074
rect 283 2057 285 2060
rect 1167 2052 1169 2066
rect 1613 2075 1615 2079
rect 1480 2042 1482 2055
rect 1488 2051 1490 2055
rect 1510 2042 1512 2055
rect 1518 2042 1520 2055
rect 1550 2054 1552 2058
rect 1573 2052 1575 2071
rect 1167 2039 1169 2042
rect 1573 2038 1575 2043
rect 1581 2038 1583 2042
rect 1613 2041 1615 2055
rect 1480 2028 1482 2032
rect 1510 2028 1512 2032
rect 1518 2028 1520 2032
rect 1613 2028 1615 2031
rect 1573 2024 1575 2028
rect 1581 2024 1583 2028
rect 150 2002 152 2006
rect 385 2005 387 2008
rect 57 1986 59 1990
rect 65 1986 67 1990
rect 87 1986 89 1990
rect 95 1986 97 1990
rect 127 1989 129 1993
rect 190 1986 192 1990
rect 57 1953 59 1966
rect 65 1962 67 1966
rect 87 1953 89 1966
rect 95 1953 97 1966
rect 127 1965 129 1969
rect 150 1963 152 1982
rect 797 2003 814 2005
rect 834 2003 847 2005
rect 867 2003 870 2005
rect 797 1995 814 1997
rect 834 1995 847 1997
rect 867 1995 870 1997
rect 273 1980 290 1982
rect 310 1980 323 1982
rect 343 1980 346 1982
rect 273 1972 290 1974
rect 310 1972 323 1974
rect 343 1972 346 1974
rect 385 1971 387 1985
rect 150 1949 152 1954
rect 158 1949 160 1953
rect 190 1952 192 1966
rect 385 1958 387 1961
rect 57 1939 59 1943
rect 87 1939 89 1943
rect 95 1939 97 1943
rect 190 1939 192 1942
rect 150 1935 152 1939
rect 158 1935 160 1939
rect 150 1861 152 1865
rect 57 1845 59 1849
rect 65 1845 67 1849
rect 87 1845 89 1849
rect 95 1845 97 1849
rect 127 1848 129 1852
rect 307 1858 309 1871
rect 330 1858 332 1862
rect 190 1845 192 1849
rect 57 1812 59 1825
rect 65 1821 67 1825
rect 87 1812 89 1825
rect 95 1812 97 1825
rect 127 1824 129 1828
rect 150 1822 152 1841
rect 698 1839 715 1841
rect 735 1839 748 1841
rect 768 1839 771 1841
rect 307 1825 309 1838
rect 330 1834 332 1838
rect 698 1831 715 1833
rect 735 1831 748 1833
rect 768 1831 771 1833
rect 1189 1827 1191 1840
rect 1212 1827 1214 1831
rect 1573 1829 1575 1833
rect 150 1808 152 1813
rect 158 1808 160 1812
rect 190 1811 192 1825
rect 283 1821 285 1824
rect 57 1798 59 1802
rect 87 1798 89 1802
rect 95 1798 97 1802
rect 330 1819 332 1826
rect 307 1812 309 1815
rect 884 1818 901 1820
rect 921 1818 934 1820
rect 964 1818 967 1820
rect 884 1810 901 1812
rect 921 1810 934 1812
rect 964 1810 967 1812
rect 330 1806 332 1809
rect 1480 1813 1482 1817
rect 1488 1813 1490 1817
rect 1510 1813 1512 1817
rect 1518 1813 1520 1817
rect 1550 1816 1552 1820
rect 884 1802 901 1804
rect 921 1802 934 1804
rect 964 1802 967 1804
rect 190 1798 192 1801
rect 150 1794 152 1798
rect 158 1794 160 1798
rect 283 1787 285 1801
rect 1189 1794 1191 1807
rect 1212 1803 1214 1807
rect 1165 1790 1167 1793
rect 283 1774 285 1777
rect 692 1773 709 1775
rect 729 1773 742 1775
rect 772 1773 775 1775
rect 1212 1788 1214 1795
rect 1613 1813 1615 1817
rect 1189 1781 1191 1784
rect 1480 1780 1482 1793
rect 1488 1789 1490 1793
rect 1510 1780 1512 1793
rect 1518 1780 1520 1793
rect 1550 1792 1552 1796
rect 1573 1790 1575 1809
rect 1212 1775 1214 1778
rect 1573 1776 1575 1781
rect 1581 1776 1583 1780
rect 1613 1779 1615 1793
rect 692 1765 709 1767
rect 729 1765 742 1767
rect 772 1765 775 1767
rect 692 1757 709 1759
rect 729 1757 742 1759
rect 772 1757 775 1759
rect 1165 1756 1167 1770
rect 1480 1766 1482 1770
rect 1510 1766 1512 1770
rect 1518 1766 1520 1770
rect 1613 1766 1615 1769
rect 1573 1762 1575 1766
rect 1581 1762 1583 1766
rect 1165 1743 1167 1746
rect 150 1719 152 1723
rect 57 1703 59 1707
rect 65 1703 67 1707
rect 87 1703 89 1707
rect 95 1703 97 1707
rect 127 1706 129 1710
rect 388 1717 390 1720
rect 190 1703 192 1707
rect 57 1670 59 1683
rect 65 1679 67 1683
rect 87 1670 89 1683
rect 95 1670 97 1683
rect 127 1682 129 1686
rect 150 1680 152 1699
rect 273 1697 290 1699
rect 310 1697 323 1699
rect 343 1697 346 1699
rect 273 1689 290 1691
rect 310 1689 323 1691
rect 343 1689 346 1691
rect 388 1683 390 1697
rect 150 1666 152 1671
rect 158 1666 160 1670
rect 190 1669 192 1683
rect 388 1670 390 1673
rect 57 1656 59 1660
rect 87 1656 89 1660
rect 95 1656 97 1660
rect 190 1656 192 1659
rect 150 1652 152 1656
rect 158 1652 160 1656
rect 706 1565 723 1567
rect 743 1565 756 1567
rect 776 1565 779 1567
rect 706 1557 723 1559
rect 743 1557 756 1559
rect 776 1557 779 1559
rect 150 1532 152 1536
rect 57 1516 59 1520
rect 65 1516 67 1520
rect 87 1516 89 1520
rect 95 1516 97 1520
rect 127 1519 129 1523
rect 307 1529 309 1542
rect 330 1529 332 1533
rect 190 1516 192 1520
rect 57 1483 59 1496
rect 65 1492 67 1496
rect 87 1483 89 1496
rect 95 1483 97 1496
rect 127 1495 129 1499
rect 150 1493 152 1512
rect 307 1496 309 1509
rect 330 1505 332 1509
rect 700 1499 717 1501
rect 737 1499 750 1501
rect 780 1499 783 1501
rect 150 1479 152 1484
rect 158 1479 160 1483
rect 190 1482 192 1496
rect 283 1492 285 1495
rect 57 1469 59 1473
rect 87 1469 89 1473
rect 95 1469 97 1473
rect 330 1490 332 1497
rect 700 1491 717 1493
rect 737 1491 750 1493
rect 780 1491 783 1493
rect 307 1483 309 1486
rect 893 1487 910 1489
rect 930 1487 943 1489
rect 983 1487 986 1489
rect 700 1483 717 1485
rect 737 1483 750 1485
rect 780 1483 783 1485
rect 330 1477 332 1480
rect 893 1479 910 1481
rect 930 1479 943 1481
rect 983 1479 986 1481
rect 190 1469 192 1472
rect 150 1465 152 1469
rect 158 1465 160 1469
rect 283 1458 285 1472
rect 893 1471 910 1473
rect 930 1471 943 1473
rect 983 1471 986 1473
rect 1189 1467 1191 1480
rect 1212 1467 1214 1471
rect 893 1463 910 1465
rect 930 1463 943 1465
rect 983 1463 986 1465
rect 283 1445 285 1448
rect 1573 1462 1575 1466
rect 1189 1434 1191 1447
rect 1212 1443 1214 1447
rect 1480 1446 1482 1450
rect 1488 1446 1490 1450
rect 1510 1446 1512 1450
rect 1518 1446 1520 1450
rect 1550 1449 1552 1453
rect 1165 1430 1167 1433
rect 700 1417 717 1419
rect 737 1417 750 1419
rect 790 1417 793 1419
rect 700 1409 717 1411
rect 737 1409 750 1411
rect 790 1409 793 1411
rect 1212 1428 1214 1435
rect 1189 1421 1191 1424
rect 1613 1446 1615 1450
rect 1212 1415 1214 1418
rect 1480 1413 1482 1426
rect 1488 1422 1490 1426
rect 1510 1413 1512 1426
rect 1518 1413 1520 1426
rect 1550 1425 1552 1429
rect 1573 1423 1575 1442
rect 700 1401 717 1403
rect 737 1401 750 1403
rect 790 1401 793 1403
rect 150 1390 152 1394
rect 388 1391 390 1394
rect 1165 1396 1167 1410
rect 1573 1409 1575 1414
rect 1581 1409 1583 1413
rect 1613 1412 1615 1426
rect 1480 1400 1482 1403
rect 1510 1399 1512 1403
rect 1518 1399 1520 1403
rect 1613 1399 1615 1402
rect 700 1393 717 1395
rect 737 1393 750 1395
rect 790 1393 793 1395
rect 57 1374 59 1378
rect 65 1374 67 1378
rect 87 1374 89 1378
rect 95 1374 97 1378
rect 127 1377 129 1381
rect 190 1374 192 1378
rect 57 1341 59 1354
rect 65 1350 67 1354
rect 87 1341 89 1354
rect 95 1341 97 1354
rect 127 1353 129 1357
rect 150 1351 152 1370
rect 1573 1395 1575 1399
rect 1581 1395 1583 1399
rect 1165 1383 1167 1386
rect 273 1368 290 1370
rect 310 1368 323 1370
rect 343 1368 346 1370
rect 273 1360 290 1362
rect 310 1360 323 1362
rect 343 1360 346 1362
rect 388 1357 390 1371
rect 150 1337 152 1342
rect 158 1337 160 1341
rect 190 1340 192 1354
rect 388 1344 390 1347
rect 57 1327 59 1331
rect 87 1327 89 1331
rect 95 1327 97 1331
rect 190 1327 192 1330
rect 150 1323 152 1327
rect 158 1323 160 1327
rect 708 1151 725 1153
rect 745 1151 758 1153
rect 778 1151 781 1153
rect 708 1143 725 1145
rect 745 1143 758 1145
rect 778 1143 781 1145
rect 702 1085 719 1087
rect 739 1085 752 1087
rect 782 1085 785 1087
rect 702 1077 719 1079
rect 739 1077 752 1079
rect 782 1077 785 1079
rect 702 1069 719 1071
rect 739 1069 752 1071
rect 782 1069 785 1071
rect 150 1042 152 1046
rect 57 1026 59 1030
rect 65 1026 67 1030
rect 87 1026 89 1030
rect 95 1026 97 1030
rect 127 1029 129 1033
rect 305 1040 307 1053
rect 1189 1052 1191 1065
rect 1212 1052 1214 1056
rect 328 1040 330 1044
rect 190 1026 192 1030
rect 57 993 59 1006
rect 65 1002 67 1006
rect 87 993 89 1006
rect 95 993 97 1006
rect 127 1005 129 1009
rect 150 1003 152 1022
rect 918 1032 941 1034
rect 955 1032 968 1034
rect 1018 1032 1021 1034
rect 1573 1044 1575 1048
rect 918 1024 941 1026
rect 955 1024 968 1026
rect 1018 1024 1021 1026
rect 305 1007 307 1020
rect 328 1016 330 1020
rect 1189 1019 1191 1032
rect 1212 1028 1214 1032
rect 1480 1028 1482 1032
rect 1488 1028 1490 1032
rect 1510 1028 1512 1032
rect 1518 1028 1520 1032
rect 1550 1031 1552 1035
rect 918 1016 941 1018
rect 955 1016 968 1018
rect 1018 1016 1021 1018
rect 150 989 152 994
rect 158 989 160 993
rect 190 992 192 1006
rect 281 1003 283 1006
rect 57 979 59 983
rect 87 979 89 983
rect 95 979 97 983
rect 328 1001 330 1008
rect 1165 1015 1167 1018
rect 918 1008 941 1010
rect 955 1008 968 1010
rect 1018 1008 1021 1010
rect 702 1003 719 1005
rect 739 1003 752 1005
rect 792 1003 795 1005
rect 305 994 307 997
rect 918 1000 941 1002
rect 955 1000 968 1002
rect 1018 1000 1021 1002
rect 702 995 719 997
rect 739 995 752 997
rect 792 995 795 997
rect 1212 1013 1214 1020
rect 1189 1006 1191 1009
rect 1613 1028 1615 1032
rect 1212 1000 1214 1003
rect 1480 995 1482 1008
rect 1488 1004 1490 1008
rect 1510 995 1512 1008
rect 1518 995 1520 1008
rect 1550 1007 1552 1011
rect 1573 1005 1575 1024
rect 328 988 330 991
rect 702 987 719 989
rect 739 987 752 989
rect 792 987 795 989
rect 190 979 192 982
rect 150 975 152 979
rect 158 975 160 979
rect 281 969 283 983
rect 1165 981 1167 995
rect 1573 991 1575 996
rect 1581 991 1583 995
rect 1613 994 1615 1008
rect 1480 981 1482 985
rect 1510 981 1512 985
rect 1518 981 1520 985
rect 1613 981 1615 984
rect 702 979 719 981
rect 739 979 752 981
rect 792 979 795 981
rect 1573 977 1575 981
rect 1581 977 1583 981
rect 1165 968 1167 971
rect 281 956 283 959
rect 703 916 726 918
rect 740 916 753 918
rect 803 916 806 918
rect 387 906 389 909
rect 703 908 726 910
rect 740 908 753 910
rect 803 908 806 910
rect 148 901 150 905
rect 55 885 57 889
rect 63 885 65 889
rect 85 885 87 889
rect 93 885 95 889
rect 125 888 127 892
rect 188 885 190 889
rect 703 900 726 902
rect 740 900 753 902
rect 803 900 806 902
rect 703 892 726 894
rect 740 892 753 894
rect 803 892 806 894
rect 55 852 57 865
rect 63 861 65 865
rect 85 852 87 865
rect 93 852 95 865
rect 125 864 127 868
rect 148 862 150 881
rect 271 879 288 881
rect 308 879 321 881
rect 341 879 344 881
rect 271 871 288 873
rect 308 871 321 873
rect 341 871 344 873
rect 387 872 389 886
rect 703 884 726 886
rect 740 884 753 886
rect 803 884 806 886
rect 148 848 150 853
rect 156 848 158 852
rect 188 851 190 865
rect 387 859 389 862
rect 55 838 57 842
rect 85 838 87 842
rect 93 838 95 842
rect 188 838 190 841
rect 148 834 150 838
rect 156 834 158 838
rect 707 656 724 658
rect 744 656 757 658
rect 777 656 780 658
rect 707 648 724 650
rect 744 648 757 650
rect 777 648 780 650
rect 701 590 718 592
rect 738 590 751 592
rect 781 590 784 592
rect 701 582 718 584
rect 738 582 751 584
rect 781 582 784 584
rect 701 574 718 576
rect 738 574 751 576
rect 781 574 784 576
rect 148 552 150 556
rect 55 536 57 540
rect 63 536 65 540
rect 85 536 87 540
rect 93 536 95 540
rect 125 539 127 543
rect 304 550 306 563
rect 327 550 329 554
rect 188 536 190 540
rect 55 503 57 516
rect 63 512 65 516
rect 85 503 87 516
rect 93 503 95 516
rect 125 515 127 519
rect 148 513 150 532
rect 304 517 306 530
rect 327 526 329 530
rect 925 524 942 526
rect 962 524 975 526
rect 1035 524 1038 526
rect 148 499 150 504
rect 156 499 158 503
rect 188 502 190 516
rect 280 513 282 516
rect 55 489 57 493
rect 85 489 87 493
rect 93 489 95 493
rect 327 511 329 518
rect 925 516 942 518
rect 962 516 975 518
rect 1035 516 1038 518
rect 304 504 306 507
rect 701 508 718 510
rect 738 508 751 510
rect 791 508 794 510
rect 1189 512 1191 525
rect 1212 512 1214 516
rect 925 508 942 510
rect 962 508 975 510
rect 1035 508 1038 510
rect 327 498 329 501
rect 701 500 718 502
rect 738 500 751 502
rect 791 500 794 502
rect 925 500 942 502
rect 962 500 975 502
rect 1035 500 1038 502
rect 188 489 190 492
rect 148 485 150 489
rect 156 485 158 489
rect 280 479 282 493
rect 701 492 718 494
rect 738 492 751 494
rect 791 492 794 494
rect 925 492 942 494
rect 962 492 975 494
rect 1035 492 1038 494
rect 701 484 718 486
rect 738 484 751 486
rect 791 484 794 486
rect 925 484 942 486
rect 962 484 975 486
rect 1035 484 1038 486
rect 1189 479 1191 492
rect 1212 488 1214 492
rect 1165 475 1167 478
rect 280 466 282 469
rect 1212 473 1214 480
rect 1189 466 1191 469
rect 1573 468 1575 472
rect 1212 460 1214 463
rect 1165 441 1167 455
rect 1480 452 1482 456
rect 1488 452 1490 456
rect 1510 452 1512 456
rect 1518 452 1520 456
rect 1550 455 1552 459
rect 1613 452 1615 456
rect 1165 428 1167 431
rect 387 420 389 423
rect 702 421 725 423
rect 739 421 752 423
rect 802 421 805 423
rect 148 411 150 415
rect 55 395 57 399
rect 63 395 65 399
rect 85 395 87 399
rect 93 395 95 399
rect 125 398 127 402
rect 1480 419 1482 432
rect 1488 428 1490 432
rect 1510 419 1512 432
rect 1518 419 1520 432
rect 1550 431 1552 435
rect 1573 429 1575 448
rect 702 413 725 415
rect 739 413 752 415
rect 802 413 805 415
rect 1573 415 1575 420
rect 1581 415 1583 419
rect 1613 418 1615 432
rect 702 405 725 407
rect 739 405 752 407
rect 802 405 805 407
rect 1480 405 1482 409
rect 1510 405 1512 409
rect 1518 405 1520 409
rect 1613 405 1615 408
rect 188 395 190 399
rect 55 362 57 375
rect 63 371 65 375
rect 85 362 87 375
rect 93 362 95 375
rect 125 374 127 378
rect 148 372 150 391
rect 270 389 287 391
rect 307 389 320 391
rect 340 389 343 391
rect 387 386 389 400
rect 1573 401 1575 405
rect 1581 401 1583 405
rect 702 397 725 399
rect 739 397 752 399
rect 802 397 805 399
rect 702 389 725 391
rect 739 389 752 391
rect 802 389 805 391
rect 270 381 287 383
rect 307 381 320 383
rect 340 381 343 383
rect 148 358 150 363
rect 156 358 158 362
rect 188 361 190 375
rect 387 373 389 376
rect 55 348 57 352
rect 85 348 87 352
rect 93 348 95 352
rect 188 348 190 351
rect 148 344 150 348
rect 156 344 158 348
rect 698 317 715 319
rect 735 317 748 319
rect 808 317 811 319
rect 698 309 715 311
rect 735 309 748 311
rect 808 309 811 311
rect 698 301 715 303
rect 735 301 748 303
rect 808 301 811 303
rect 698 293 715 295
rect 735 293 748 295
rect 808 293 811 295
rect 698 285 715 287
rect 735 285 748 287
rect 808 285 811 287
rect 698 277 715 279
rect 735 277 748 279
rect 808 277 811 279
rect 1573 178 1575 182
rect 1480 162 1482 166
rect 1488 162 1490 166
rect 1510 162 1512 166
rect 1518 162 1520 166
rect 1550 165 1552 169
rect 1613 162 1615 166
rect 1480 129 1482 142
rect 1488 138 1490 142
rect 1510 129 1512 142
rect 1518 129 1520 142
rect 1550 141 1552 145
rect 1573 139 1575 158
rect 1573 125 1575 130
rect 1581 125 1583 129
rect 1613 128 1615 142
rect 1480 115 1482 119
rect 1510 115 1512 119
rect 1518 115 1520 119
rect 1613 115 1615 118
rect 1573 111 1575 115
rect 1581 111 1583 115
rect 148 82 150 86
rect 55 66 57 70
rect 63 66 65 70
rect 85 66 87 70
rect 93 66 95 70
rect 125 69 127 73
rect 188 66 190 70
rect 55 33 57 46
rect 63 42 65 46
rect 85 33 87 46
rect 93 33 95 46
rect 125 45 127 49
rect 148 43 150 62
rect 148 29 150 34
rect 156 29 158 33
rect 188 32 190 46
rect 55 19 57 23
rect 85 19 87 23
rect 93 19 95 23
rect 188 19 190 22
rect 148 15 150 19
rect 156 15 158 19
<< polycontact >>
rect 307 2154 311 2158
rect 327 2145 332 2150
rect 59 2128 63 2132
rect 96 2128 100 2132
rect 129 2131 133 2135
rect 148 2113 152 2117
rect 148 2101 152 2105
rect 1191 2136 1195 2140
rect 1211 2127 1216 2132
rect 148 2090 152 2094
rect 188 2093 192 2097
rect 697 2100 701 2104
rect 697 2092 701 2096
rect 330 2085 334 2089
rect 279 2073 283 2077
rect 1517 2079 1521 2083
rect 1550 2082 1554 2086
rect 1214 2067 1218 2071
rect 1163 2055 1167 2059
rect 1569 2064 1573 2068
rect 1476 2046 1480 2050
rect 1569 2052 1573 2056
rect 1569 2041 1573 2045
rect 1609 2044 1613 2048
rect 57 1990 61 1994
rect 94 1990 98 1994
rect 127 1993 131 1997
rect 146 1975 150 1979
rect 146 1963 150 1967
rect 269 1980 273 1984
rect 793 2003 797 2007
rect 793 1995 797 1999
rect 269 1972 273 1976
rect 381 1974 385 1978
rect 146 1952 150 1956
rect 186 1955 190 1959
rect 307 1871 311 1875
rect 57 1849 61 1853
rect 94 1849 98 1853
rect 127 1852 131 1856
rect 327 1862 332 1867
rect 146 1834 150 1838
rect 146 1822 150 1826
rect 694 1839 698 1843
rect 1189 1840 1193 1844
rect 694 1831 698 1835
rect 1209 1831 1214 1836
rect 146 1811 150 1815
rect 186 1814 190 1818
rect 880 1818 884 1822
rect 880 1810 884 1814
rect 330 1802 334 1806
rect 880 1802 884 1806
rect 1517 1817 1521 1821
rect 1550 1820 1554 1824
rect 279 1790 283 1794
rect 688 1773 692 1777
rect 688 1765 692 1769
rect 1569 1802 1573 1806
rect 1475 1784 1480 1789
rect 1569 1790 1573 1794
rect 1212 1771 1216 1775
rect 1569 1779 1573 1783
rect 1609 1782 1613 1786
rect 688 1757 692 1761
rect 1161 1759 1165 1763
rect 57 1707 61 1711
rect 94 1707 98 1711
rect 127 1710 131 1714
rect 146 1692 150 1696
rect 146 1680 150 1684
rect 269 1697 273 1701
rect 269 1689 273 1693
rect 384 1686 388 1690
rect 146 1669 150 1673
rect 186 1672 190 1676
rect 702 1565 706 1569
rect 702 1557 706 1561
rect 307 1542 311 1546
rect 57 1520 61 1524
rect 94 1520 98 1524
rect 127 1523 131 1527
rect 327 1533 332 1538
rect 146 1505 150 1509
rect 146 1493 150 1497
rect 696 1499 700 1503
rect 146 1482 150 1486
rect 186 1485 190 1489
rect 696 1491 700 1495
rect 696 1483 700 1487
rect 889 1487 893 1491
rect 889 1479 893 1483
rect 1189 1480 1193 1484
rect 330 1473 334 1477
rect 279 1461 283 1465
rect 889 1471 893 1475
rect 889 1463 893 1467
rect 1209 1471 1214 1476
rect 1517 1450 1521 1454
rect 1550 1453 1554 1457
rect 696 1417 700 1421
rect 696 1409 700 1413
rect 1569 1435 1573 1439
rect 1475 1417 1480 1422
rect 1212 1411 1216 1415
rect 1569 1423 1573 1427
rect 696 1401 700 1405
rect 696 1393 700 1397
rect 1161 1399 1165 1403
rect 1569 1412 1573 1416
rect 1609 1415 1613 1419
rect 57 1378 61 1382
rect 94 1378 98 1382
rect 127 1381 131 1385
rect 146 1363 150 1367
rect 146 1351 150 1355
rect 269 1368 273 1372
rect 269 1360 273 1364
rect 384 1360 388 1364
rect 146 1340 150 1344
rect 186 1343 190 1347
rect 704 1151 708 1155
rect 704 1143 708 1147
rect 698 1085 702 1089
rect 698 1077 702 1081
rect 698 1069 702 1073
rect 1189 1065 1193 1069
rect 305 1053 309 1057
rect 57 1030 61 1034
rect 94 1030 98 1034
rect 127 1033 131 1037
rect 1209 1056 1214 1061
rect 325 1044 330 1049
rect 146 1015 150 1019
rect 146 1003 150 1007
rect 914 1031 918 1035
rect 1517 1032 1521 1036
rect 1550 1035 1554 1039
rect 914 1023 918 1027
rect 914 1015 918 1019
rect 146 992 150 996
rect 186 995 190 999
rect 698 1003 702 1007
rect 914 1007 918 1011
rect 698 995 702 999
rect 914 999 918 1003
rect 1569 1017 1573 1021
rect 1212 996 1216 1000
rect 1475 999 1480 1004
rect 1569 1005 1573 1009
rect 328 984 332 988
rect 698 987 702 991
rect 277 972 281 976
rect 698 979 702 983
rect 1161 984 1165 988
rect 1569 994 1573 998
rect 1609 997 1613 1001
rect 699 915 703 919
rect 699 907 703 911
rect 55 889 59 893
rect 92 889 96 893
rect 125 892 129 896
rect 699 899 703 903
rect 699 891 703 895
rect 144 874 148 878
rect 144 862 148 866
rect 267 879 271 883
rect 267 871 271 875
rect 383 875 387 879
rect 699 881 703 886
rect 144 851 148 855
rect 184 854 188 858
rect 703 656 707 660
rect 703 648 707 652
rect 697 590 701 594
rect 697 582 701 586
rect 697 574 701 578
rect 304 563 308 567
rect 55 540 59 544
rect 92 540 96 544
rect 125 543 129 547
rect 324 554 329 559
rect 144 525 148 529
rect 144 513 148 517
rect 921 524 925 528
rect 1189 525 1193 529
rect 144 502 148 506
rect 184 505 188 509
rect 921 516 925 520
rect 697 508 701 512
rect 921 508 925 512
rect 1209 516 1214 521
rect 697 500 701 504
rect 921 500 925 504
rect 327 494 331 498
rect 276 482 280 486
rect 697 492 701 496
rect 921 492 925 496
rect 697 484 701 488
rect 921 484 925 488
rect 1212 456 1216 460
rect 1517 456 1521 460
rect 1550 459 1554 463
rect 1161 444 1165 448
rect 1569 441 1573 445
rect 698 420 702 424
rect 1475 423 1480 428
rect 55 399 59 403
rect 92 399 96 403
rect 125 402 129 406
rect 698 412 702 416
rect 1569 429 1573 433
rect 698 404 702 408
rect 1569 418 1573 422
rect 1609 421 1613 425
rect 144 384 148 388
rect 144 372 148 376
rect 266 389 270 393
rect 383 389 387 393
rect 266 381 270 385
rect 698 396 702 400
rect 698 387 702 391
rect 144 361 148 365
rect 184 364 188 368
rect 694 317 698 321
rect 694 309 698 313
rect 694 301 698 305
rect 694 293 698 297
rect 694 284 698 288
rect 694 275 698 279
rect 1480 166 1484 170
rect 1517 166 1521 170
rect 1550 169 1554 173
rect 1569 151 1573 155
rect 1475 133 1480 138
rect 1569 139 1573 143
rect 1569 128 1573 132
rect 1609 131 1613 135
rect 55 70 59 74
rect 92 70 96 74
rect 125 73 129 77
rect 144 55 148 59
rect 144 43 148 47
rect 144 32 148 36
rect 184 35 188 39
<< metal1 >>
rect 25 2186 565 2189
rect 25 2058 28 2186
rect 249 2166 311 2170
rect 51 2148 197 2152
rect 201 2148 204 2152
rect 51 2120 54 2148
rect 59 2132 63 2135
rect 81 2120 84 2148
rect 92 2140 103 2145
rect 96 2132 101 2140
rect 100 2128 101 2132
rect 121 2120 124 2148
rect 147 2140 151 2148
rect 129 2135 133 2138
rect 136 2124 142 2127
rect 139 2117 142 2124
rect 139 2113 148 2117
rect 70 2101 74 2104
rect 100 2100 104 2104
rect 143 2101 148 2105
rect 143 2100 147 2101
rect 100 2096 147 2100
rect 70 2091 74 2096
rect 100 2091 104 2096
rect 143 2094 147 2096
rect 163 2097 167 2120
rect 187 2124 191 2148
rect 195 2097 199 2104
rect 249 2097 253 2166
rect 307 2159 311 2166
rect 307 2158 350 2159
rect 311 2154 350 2158
rect 302 2145 327 2150
rect 267 2141 306 2145
rect 267 2128 271 2141
rect 268 2121 271 2128
rect 143 2090 148 2094
rect 163 2093 188 2097
rect 195 2093 253 2097
rect 163 2087 167 2093
rect 195 2090 199 2093
rect 54 2063 58 2081
rect 84 2063 89 2081
rect 147 2063 151 2077
rect 187 2063 191 2080
rect 267 2077 271 2121
rect 279 2112 283 2117
rect 310 2115 314 2121
rect 325 2115 329 2121
rect 310 2111 329 2115
rect 310 2108 314 2111
rect 278 2104 282 2108
rect 286 2077 290 2084
rect 317 2104 321 2111
rect 325 2102 329 2111
rect 302 2077 306 2098
rect 333 2115 337 2121
rect 345 2115 350 2154
rect 333 2111 350 2115
rect 333 2102 337 2111
rect 433 2095 437 2157
rect 441 2106 445 2162
rect 330 2077 334 2085
rect 267 2073 279 2077
rect 286 2073 334 2077
rect 286 2070 290 2073
rect 38 2058 42 2063
rect 46 2058 266 2063
rect 23 2052 44 2058
rect 261 2057 266 2058
rect 278 2057 282 2060
rect 261 2056 282 2057
rect 261 2052 278 2056
rect 38 1925 44 2052
rect 49 2010 195 2014
rect 199 2010 202 2014
rect 49 1982 52 2010
rect 57 1994 61 1997
rect 79 1982 82 2010
rect 90 2002 101 2007
rect 94 1994 99 2002
rect 98 1990 99 1994
rect 119 1982 122 2010
rect 145 2002 149 2010
rect 134 1986 140 1989
rect 137 1979 140 1986
rect 137 1975 146 1979
rect 68 1963 72 1966
rect 98 1962 102 1966
rect 141 1963 146 1967
rect 141 1962 145 1963
rect 98 1958 145 1962
rect 68 1953 72 1958
rect 98 1953 102 1958
rect 141 1956 145 1958
rect 161 1959 165 1982
rect 185 1986 189 2010
rect 380 2005 384 2009
rect 316 1992 367 1996
rect 316 1987 320 1992
rect 193 1959 197 1966
rect 281 1983 290 1987
rect 316 1983 323 1987
rect 210 1972 269 1976
rect 210 1959 214 1972
rect 281 1971 285 1983
rect 316 1979 320 1983
rect 310 1975 320 1979
rect 363 1978 367 1992
rect 388 1978 392 1985
rect 363 1974 381 1978
rect 388 1974 398 1978
rect 285 1967 290 1971
rect 343 1967 347 1971
rect 388 1971 392 1974
rect 141 1952 146 1956
rect 161 1955 186 1959
rect 193 1955 214 1959
rect 161 1949 165 1955
rect 193 1952 197 1955
rect 52 1925 56 1943
rect 82 1925 87 1943
rect 145 1925 149 1939
rect 185 1925 189 1942
rect 347 1925 351 1967
rect 380 1957 384 1961
rect 380 1925 384 1953
rect 38 1920 40 1925
rect 44 1920 384 1925
rect 38 1784 44 1920
rect 251 1881 311 1885
rect 49 1869 195 1873
rect 199 1869 202 1873
rect 49 1841 52 1869
rect 57 1853 61 1856
rect 79 1841 82 1869
rect 90 1861 101 1866
rect 94 1853 99 1861
rect 98 1849 99 1853
rect 119 1841 122 1869
rect 145 1861 149 1869
rect 134 1845 140 1848
rect 137 1838 140 1845
rect 137 1834 146 1838
rect 68 1822 72 1825
rect 98 1821 102 1825
rect 141 1822 146 1826
rect 141 1821 145 1822
rect 98 1817 145 1821
rect 68 1812 72 1817
rect 98 1812 102 1817
rect 141 1815 145 1817
rect 161 1818 165 1841
rect 185 1845 189 1869
rect 193 1818 197 1825
rect 251 1819 255 1881
rect 307 1876 311 1881
rect 307 1875 350 1876
rect 311 1871 350 1875
rect 302 1862 327 1867
rect 267 1858 306 1862
rect 141 1811 146 1815
rect 161 1814 186 1818
rect 193 1814 251 1818
rect 161 1808 165 1814
rect 193 1811 197 1814
rect 52 1784 56 1802
rect 82 1784 87 1802
rect 145 1784 149 1798
rect 185 1784 189 1801
rect 267 1794 271 1858
rect 279 1829 283 1834
rect 310 1832 314 1838
rect 325 1832 329 1838
rect 310 1828 329 1832
rect 310 1825 314 1828
rect 278 1821 282 1825
rect 286 1794 290 1801
rect 317 1821 321 1828
rect 325 1819 329 1828
rect 302 1794 306 1815
rect 333 1832 337 1838
rect 345 1832 350 1871
rect 333 1828 350 1832
rect 333 1819 337 1828
rect 330 1794 334 1802
rect 267 1790 279 1794
rect 286 1790 334 1794
rect 286 1787 290 1790
rect 38 1779 40 1784
rect 44 1779 258 1784
rect 38 1642 44 1779
rect 253 1774 258 1779
rect 278 1774 282 1777
rect 253 1773 282 1774
rect 253 1769 278 1773
rect 433 1761 437 2090
rect 441 2069 445 2101
rect 441 1770 445 2064
rect 449 1978 453 2162
rect 449 1834 453 1973
rect 457 1999 461 2162
rect 457 1969 461 1994
rect 49 1727 195 1731
rect 199 1727 202 1731
rect 49 1699 52 1727
rect 57 1711 61 1714
rect 79 1699 82 1727
rect 90 1719 101 1724
rect 94 1711 99 1719
rect 98 1707 99 1711
rect 119 1699 122 1727
rect 145 1719 149 1727
rect 134 1703 140 1706
rect 137 1696 140 1703
rect 137 1692 146 1696
rect 68 1680 72 1683
rect 98 1679 102 1683
rect 141 1680 146 1684
rect 141 1679 145 1680
rect 98 1675 145 1679
rect 68 1670 72 1675
rect 98 1670 102 1675
rect 141 1673 145 1675
rect 161 1676 165 1699
rect 185 1703 189 1727
rect 383 1717 387 1721
rect 316 1713 368 1717
rect 316 1704 320 1713
rect 267 1697 269 1701
rect 281 1700 290 1704
rect 316 1700 323 1704
rect 193 1676 197 1683
rect 222 1690 269 1693
rect 217 1689 269 1690
rect 217 1676 221 1689
rect 281 1688 285 1700
rect 316 1696 320 1700
rect 310 1692 320 1696
rect 364 1690 368 1713
rect 391 1690 395 1697
rect 285 1684 290 1688
rect 343 1684 347 1688
rect 364 1686 384 1690
rect 391 1686 405 1690
rect 141 1669 146 1673
rect 161 1672 186 1676
rect 193 1672 221 1676
rect 161 1666 165 1672
rect 193 1669 197 1672
rect 52 1642 56 1660
rect 82 1642 87 1660
rect 145 1642 149 1656
rect 185 1642 189 1659
rect 347 1642 352 1684
rect 391 1683 395 1686
rect 383 1669 387 1673
rect 382 1642 387 1665
rect 38 1637 40 1642
rect 44 1637 387 1642
rect 38 1455 44 1637
rect 249 1553 311 1557
rect 49 1540 195 1544
rect 199 1540 202 1544
rect 49 1512 52 1540
rect 57 1524 61 1527
rect 79 1512 82 1540
rect 90 1532 101 1537
rect 94 1524 99 1532
rect 98 1520 99 1524
rect 119 1512 122 1540
rect 145 1532 149 1540
rect 134 1516 140 1519
rect 137 1509 140 1516
rect 137 1505 146 1509
rect 68 1493 72 1496
rect 98 1492 102 1496
rect 141 1493 146 1497
rect 141 1492 145 1493
rect 98 1488 145 1492
rect 68 1483 72 1488
rect 98 1483 102 1488
rect 141 1486 145 1488
rect 161 1489 165 1512
rect 185 1516 189 1540
rect 193 1489 197 1496
rect 249 1490 253 1553
rect 307 1547 311 1553
rect 307 1546 350 1547
rect 311 1542 350 1546
rect 302 1533 327 1538
rect 267 1529 306 1533
rect 141 1482 146 1486
rect 161 1485 186 1489
rect 193 1485 249 1489
rect 161 1479 165 1485
rect 193 1482 197 1485
rect 52 1455 56 1473
rect 82 1455 87 1473
rect 145 1455 149 1469
rect 185 1455 189 1472
rect 267 1465 271 1529
rect 279 1500 283 1505
rect 310 1503 314 1509
rect 325 1503 329 1509
rect 310 1499 329 1503
rect 310 1496 314 1499
rect 278 1492 282 1496
rect 286 1465 290 1472
rect 317 1492 321 1499
rect 325 1490 329 1499
rect 302 1465 306 1486
rect 333 1503 337 1509
rect 345 1503 350 1542
rect 333 1499 350 1503
rect 333 1490 337 1499
rect 330 1465 334 1473
rect 267 1461 279 1465
rect 286 1461 334 1465
rect 286 1458 290 1461
rect 38 1450 40 1455
rect 44 1450 257 1455
rect 38 1313 44 1450
rect 252 1445 257 1450
rect 278 1445 282 1448
rect 252 1444 282 1445
rect 252 1440 278 1444
rect 49 1398 195 1402
rect 199 1398 202 1402
rect 49 1370 52 1398
rect 57 1382 61 1385
rect 79 1370 82 1398
rect 90 1390 101 1395
rect 94 1382 99 1390
rect 98 1378 99 1382
rect 119 1370 122 1398
rect 145 1390 149 1398
rect 134 1374 140 1377
rect 137 1367 140 1374
rect 137 1363 146 1367
rect 68 1351 72 1354
rect 98 1350 102 1354
rect 141 1351 146 1355
rect 141 1350 145 1351
rect 98 1346 145 1350
rect 68 1341 72 1346
rect 98 1341 102 1346
rect 141 1344 145 1346
rect 161 1347 165 1370
rect 185 1374 189 1398
rect 383 1391 387 1395
rect 433 1395 437 1756
rect 441 1404 445 1765
rect 449 1486 453 1829
rect 316 1384 367 1388
rect 316 1375 320 1384
rect 268 1368 269 1372
rect 281 1371 290 1375
rect 316 1371 323 1375
rect 193 1347 197 1354
rect 250 1360 269 1364
rect 141 1340 146 1344
rect 161 1343 186 1347
rect 193 1343 212 1347
rect 250 1347 254 1360
rect 281 1359 285 1371
rect 316 1367 320 1371
rect 310 1363 320 1367
rect 363 1364 367 1384
rect 391 1364 395 1371
rect 363 1360 384 1364
rect 391 1360 405 1364
rect 285 1355 290 1359
rect 343 1355 347 1359
rect 391 1357 395 1360
rect 219 1343 254 1347
rect 161 1337 165 1343
rect 193 1340 197 1343
rect 52 1313 56 1331
rect 82 1313 87 1331
rect 145 1313 149 1327
rect 185 1313 189 1330
rect 347 1313 352 1355
rect 383 1343 387 1347
rect 382 1313 387 1339
rect 38 1308 40 1313
rect 44 1308 387 1313
rect 38 965 44 1308
rect 250 1063 309 1067
rect 49 1050 195 1054
rect 199 1050 202 1054
rect 49 1022 52 1050
rect 57 1034 61 1037
rect 79 1022 82 1050
rect 90 1042 101 1047
rect 94 1034 99 1042
rect 98 1030 99 1034
rect 119 1022 122 1050
rect 145 1042 149 1050
rect 134 1026 140 1029
rect 137 1019 140 1026
rect 137 1015 146 1019
rect 68 1003 72 1006
rect 98 1002 102 1006
rect 141 1003 146 1007
rect 141 1002 145 1003
rect 98 998 145 1002
rect 68 993 72 998
rect 98 993 102 998
rect 141 996 145 998
rect 161 999 165 1022
rect 185 1026 189 1050
rect 193 999 197 1006
rect 250 999 254 1063
rect 305 1058 309 1063
rect 305 1057 348 1058
rect 309 1053 348 1057
rect 300 1044 325 1049
rect 265 1040 304 1044
rect 265 1016 269 1040
rect 265 1011 271 1016
rect 279 1011 283 1016
rect 308 1014 312 1020
rect 323 1014 327 1020
rect 141 992 146 996
rect 161 995 186 999
rect 193 995 250 999
rect 161 989 165 995
rect 193 992 197 995
rect 52 965 56 983
rect 82 965 87 983
rect 145 965 149 979
rect 185 965 189 982
rect 265 976 269 1011
rect 308 1010 327 1014
rect 308 1007 312 1010
rect 276 1003 280 1007
rect 284 976 288 983
rect 315 1003 319 1010
rect 323 1001 327 1010
rect 300 976 304 997
rect 331 1014 335 1020
rect 343 1014 348 1053
rect 331 1010 348 1014
rect 331 1001 335 1010
rect 328 976 332 984
rect 265 972 277 976
rect 284 972 332 976
rect 284 969 288 972
rect 38 960 40 965
rect 44 960 251 965
rect 38 824 44 960
rect 246 956 251 960
rect 276 956 280 959
rect 246 955 280 956
rect 246 951 276 955
rect 47 909 193 913
rect 197 909 200 913
rect 47 881 50 909
rect 55 893 59 896
rect 77 881 80 909
rect 88 901 99 906
rect 92 893 97 901
rect 96 889 97 893
rect 117 881 120 909
rect 143 901 147 909
rect 132 885 138 888
rect 135 878 138 885
rect 135 874 144 878
rect 66 862 70 865
rect 96 861 100 865
rect 139 862 144 866
rect 139 861 143 862
rect 96 857 143 861
rect 66 852 70 857
rect 96 852 100 857
rect 139 855 143 857
rect 159 858 163 881
rect 183 885 187 909
rect 382 906 386 910
rect 433 906 437 1390
rect 314 895 359 899
rect 314 886 318 895
rect 260 879 267 883
rect 279 882 288 886
rect 314 882 321 886
rect 191 858 195 865
rect 220 871 267 875
rect 215 858 219 871
rect 279 870 283 882
rect 314 878 318 882
rect 355 879 359 895
rect 390 879 394 886
rect 308 874 318 878
rect 355 875 383 879
rect 390 875 404 879
rect 390 872 394 875
rect 283 866 288 870
rect 341 866 345 870
rect 139 851 144 855
rect 159 854 184 858
rect 191 854 219 858
rect 159 848 163 854
rect 191 851 195 854
rect 50 824 54 842
rect 80 824 85 842
rect 143 824 147 838
rect 183 824 187 841
rect 344 824 349 866
rect 382 858 386 862
rect 381 824 386 854
rect 42 819 386 824
rect 38 680 44 819
rect 33 676 44 680
rect 38 475 44 676
rect 238 577 308 581
rect 47 560 193 564
rect 197 560 200 564
rect 47 532 50 560
rect 55 544 59 547
rect 77 532 80 560
rect 88 552 99 557
rect 92 544 97 552
rect 96 540 97 544
rect 117 532 120 560
rect 143 552 147 560
rect 125 547 130 552
rect 132 536 138 539
rect 135 529 138 536
rect 135 525 144 529
rect 66 513 70 516
rect 96 512 100 516
rect 139 513 144 517
rect 139 512 143 513
rect 96 508 143 512
rect 66 503 70 508
rect 96 503 100 508
rect 139 506 143 508
rect 159 509 163 532
rect 183 536 187 560
rect 191 509 195 516
rect 238 509 242 577
rect 304 568 308 577
rect 304 567 347 568
rect 308 563 347 567
rect 299 554 324 559
rect 264 550 303 554
rect 264 542 268 550
rect 265 536 268 542
rect 264 526 268 536
rect 264 521 271 526
rect 279 521 283 526
rect 307 524 311 530
rect 322 524 326 530
rect 139 502 144 506
rect 159 505 184 509
rect 191 505 238 509
rect 159 499 163 505
rect 191 502 195 505
rect 50 475 54 493
rect 80 475 85 493
rect 143 475 147 489
rect 183 475 187 492
rect 264 486 268 521
rect 307 520 326 524
rect 307 517 311 520
rect 275 513 279 517
rect 283 486 287 493
rect 314 513 318 520
rect 322 511 326 520
rect 299 486 303 507
rect 330 524 334 530
rect 342 524 347 563
rect 330 520 347 524
rect 330 511 334 520
rect 327 486 331 494
rect 264 482 276 486
rect 283 482 331 486
rect 283 479 287 482
rect 42 470 247 475
rect 38 334 44 470
rect 242 466 247 470
rect 275 466 279 469
rect 242 465 279 466
rect 242 461 275 465
rect 47 419 193 423
rect 197 419 200 423
rect 382 420 386 424
rect 47 391 50 419
rect 55 403 59 406
rect 77 391 80 419
rect 88 411 99 416
rect 92 403 97 411
rect 96 399 97 403
rect 117 391 120 419
rect 143 411 147 419
rect 132 395 138 398
rect 135 388 138 395
rect 135 384 144 388
rect 66 372 70 375
rect 96 371 100 375
rect 139 372 144 376
rect 139 371 143 372
rect 96 367 143 371
rect 66 362 70 367
rect 96 362 100 367
rect 139 365 143 367
rect 159 368 163 391
rect 183 395 187 419
rect 313 408 368 412
rect 313 396 317 408
rect 264 389 266 393
rect 278 392 287 396
rect 313 392 320 396
rect 364 393 368 408
rect 390 393 394 400
rect 191 368 195 375
rect 223 381 266 385
rect 218 368 222 381
rect 278 380 282 392
rect 313 388 317 392
rect 364 389 383 393
rect 390 389 404 393
rect 307 384 317 388
rect 390 386 394 389
rect 282 376 287 380
rect 340 376 344 380
rect 139 361 144 365
rect 159 364 184 368
rect 191 364 222 368
rect 159 358 163 364
rect 191 361 195 364
rect 50 334 54 352
rect 80 334 85 352
rect 143 334 147 348
rect 183 334 187 351
rect 344 334 349 376
rect 382 372 386 376
rect 381 334 386 368
rect 42 329 386 334
rect 38 5 44 329
rect 433 272 437 900
rect 441 893 445 1399
rect 449 981 453 1481
rect 441 288 445 888
rect 449 400 453 976
rect 47 90 193 94
rect 197 90 200 94
rect 47 62 50 90
rect 55 74 59 77
rect 77 62 80 90
rect 88 82 99 87
rect 92 74 97 82
rect 96 70 97 74
rect 117 62 120 90
rect 143 82 147 90
rect 132 66 138 69
rect 135 59 138 66
rect 135 55 144 59
rect 66 43 70 46
rect 96 42 100 46
rect 139 43 144 47
rect 139 42 143 43
rect 96 38 143 42
rect 66 33 70 38
rect 96 33 100 38
rect 139 36 143 38
rect 159 39 163 62
rect 183 66 187 90
rect 191 39 195 46
rect 433 39 437 267
rect 139 32 144 36
rect 159 35 184 39
rect 191 35 202 39
rect 159 29 163 35
rect 191 32 195 35
rect 50 5 54 23
rect 80 5 85 23
rect 143 5 147 19
rect 183 5 187 22
rect 433 16 437 34
rect 441 16 445 283
rect 449 16 453 394
rect 457 16 461 1964
rect 465 1845 469 2162
rect 465 1787 469 1840
rect 465 1778 469 1782
rect 465 1495 469 1773
rect 473 1690 477 2162
rect 473 1559 477 1685
rect 481 1801 485 2162
rect 481 1679 485 1795
rect 465 1413 469 1490
rect 465 991 469 1408
rect 473 1073 477 1554
rect 465 902 469 985
rect 465 398 469 897
rect 473 490 477 1067
rect 465 289 469 393
rect 465 16 469 284
rect 473 16 477 485
rect 481 16 485 1674
rect 489 1569 493 2162
rect 489 1504 493 1564
rect 489 1458 493 1499
rect 489 1422 493 1453
rect 489 1081 493 1417
rect 497 1364 501 2162
rect 497 1147 501 1359
rect 505 1454 509 2162
rect 505 1354 509 1449
rect 489 1013 493 1076
rect 489 911 493 1008
rect 489 495 493 906
rect 497 577 501 1142
rect 489 407 493 490
rect 489 298 493 402
rect 489 16 493 293
rect 497 16 501 572
rect 505 16 509 1349
rect 513 1156 517 2162
rect 513 1090 517 1151
rect 513 1026 517 1085
rect 513 1002 517 1020
rect 513 920 517 997
rect 513 586 517 915
rect 521 879 525 2162
rect 521 651 525 874
rect 529 1038 533 2162
rect 529 816 533 1032
rect 513 504 517 581
rect 513 416 517 499
rect 513 307 517 411
rect 513 16 517 302
rect 521 16 525 646
rect 529 16 533 811
rect 537 660 541 2162
rect 537 595 541 655
rect 537 513 541 590
rect 537 478 541 508
rect 537 425 541 473
rect 537 316 541 420
rect 545 384 549 2162
rect 537 16 541 311
rect 545 16 549 379
rect 553 543 557 2162
rect 553 325 557 538
rect 553 16 557 320
rect 561 16 565 2186
rect 1191 2140 1234 2141
rect 1195 2136 1234 2140
rect 1186 2127 1211 2132
rect 1151 2123 1190 2127
rect 744 2117 786 2121
rect 744 2107 748 2117
rect 696 2100 697 2104
rect 709 2103 718 2107
rect 744 2103 751 2107
rect 696 2092 697 2096
rect 709 2091 713 2103
rect 744 2099 748 2103
rect 738 2095 748 2099
rect 713 2087 718 2091
rect 771 2087 775 2091
rect 782 2007 786 2117
rect 1151 2059 1155 2123
rect 1194 2097 1198 2103
rect 1209 2097 1213 2103
rect 1194 2093 1213 2097
rect 1194 2090 1198 2093
rect 1162 2086 1166 2090
rect 1170 2059 1174 2066
rect 1186 2059 1190 2080
rect 1201 2072 1205 2093
rect 1209 2084 1213 2093
rect 1217 2097 1221 2103
rect 1229 2097 1234 2136
rect 1217 2093 1234 2097
rect 1217 2084 1221 2093
rect 1303 2089 1309 2210
rect 1214 2059 1218 2067
rect 1151 2055 1163 2059
rect 1170 2055 1218 2059
rect 1170 2052 1174 2055
rect 1162 2039 1166 2042
rect 840 2025 1049 2029
rect 840 2010 844 2025
rect 782 2003 793 2007
rect 805 2006 814 2010
rect 840 2006 847 2010
rect 791 1995 793 1999
rect 805 1994 809 2006
rect 840 2002 844 2006
rect 834 1998 844 2002
rect 809 1990 814 1994
rect 867 1990 870 1994
rect 1045 1880 1049 2025
rect 1045 1876 1194 1880
rect 741 1851 872 1855
rect 741 1846 745 1851
rect 692 1839 694 1843
rect 706 1842 715 1846
rect 741 1842 748 1846
rect 692 1831 694 1835
rect 706 1830 710 1842
rect 741 1838 745 1842
rect 735 1834 745 1838
rect 710 1826 715 1830
rect 768 1826 771 1830
rect 868 1822 872 1851
rect 1190 1845 1194 1876
rect 1189 1844 1232 1845
rect 1193 1840 1232 1844
rect 927 1830 1006 1834
rect 1184 1831 1209 1836
rect 927 1825 931 1830
rect 868 1818 880 1822
rect 921 1821 934 1825
rect 864 1810 880 1814
rect 892 1813 901 1817
rect 868 1802 880 1806
rect 868 1789 872 1802
rect 892 1801 896 1813
rect 927 1809 931 1821
rect 921 1805 931 1809
rect 896 1797 901 1801
rect 964 1797 967 1801
rect 735 1785 872 1789
rect 735 1780 739 1785
rect 686 1773 688 1777
rect 729 1776 742 1780
rect 686 1765 688 1769
rect 700 1768 709 1772
rect 686 1757 688 1761
rect 700 1756 704 1768
rect 735 1764 739 1776
rect 729 1760 739 1764
rect 704 1752 709 1756
rect 772 1752 775 1756
rect 749 1577 875 1581
rect 749 1572 753 1577
rect 700 1565 702 1569
rect 714 1568 723 1572
rect 749 1568 756 1572
rect 700 1557 702 1561
rect 714 1556 718 1568
rect 749 1564 753 1568
rect 743 1560 753 1564
rect 718 1552 723 1556
rect 776 1552 779 1556
rect 743 1516 853 1520
rect 743 1506 747 1516
rect 694 1499 696 1503
rect 737 1502 750 1506
rect 694 1491 696 1495
rect 708 1494 717 1498
rect 694 1483 696 1487
rect 708 1482 712 1494
rect 743 1490 747 1502
rect 737 1486 747 1490
rect 849 1483 853 1516
rect 871 1491 875 1577
rect 1002 1556 1006 1830
rect 1149 1827 1188 1831
rect 1149 1763 1153 1827
rect 1192 1801 1196 1807
rect 1207 1801 1211 1807
rect 1192 1797 1211 1801
rect 1192 1794 1196 1797
rect 1160 1790 1164 1794
rect 1168 1763 1172 1770
rect 1184 1763 1188 1784
rect 1199 1777 1203 1797
rect 1207 1788 1211 1797
rect 1215 1801 1219 1807
rect 1227 1801 1232 1840
rect 1215 1797 1232 1801
rect 1303 1822 1309 2082
rect 1338 2103 1343 2211
rect 1338 2099 1618 2103
rect 1622 2099 1626 2103
rect 1215 1788 1219 1797
rect 1212 1763 1216 1771
rect 1149 1759 1161 1763
rect 1168 1759 1216 1763
rect 1168 1756 1172 1759
rect 1160 1742 1164 1746
rect 1002 1552 1194 1556
rect 936 1500 1045 1504
rect 936 1494 940 1500
rect 871 1487 889 1491
rect 901 1490 910 1494
rect 936 1490 943 1494
rect 712 1478 717 1482
rect 780 1478 783 1482
rect 849 1479 889 1483
rect 901 1478 905 1490
rect 936 1486 940 1490
rect 930 1482 940 1486
rect 849 1471 889 1475
rect 901 1474 910 1478
rect 849 1454 853 1471
rect 871 1463 889 1467
rect 871 1434 875 1463
rect 901 1462 905 1474
rect 936 1470 940 1482
rect 930 1466 940 1470
rect 905 1458 910 1462
rect 983 1458 986 1462
rect 743 1430 875 1434
rect 743 1424 747 1430
rect 694 1417 696 1421
rect 708 1420 717 1424
rect 743 1420 750 1424
rect 694 1409 696 1413
rect 708 1408 712 1420
rect 743 1416 747 1420
rect 737 1412 747 1416
rect 694 1401 696 1405
rect 708 1404 717 1408
rect 694 1393 696 1397
rect 708 1392 712 1404
rect 743 1400 747 1412
rect 737 1396 747 1400
rect 712 1388 717 1392
rect 790 1388 793 1392
rect 751 1163 900 1167
rect 751 1158 755 1163
rect 702 1151 704 1155
rect 716 1154 725 1158
rect 751 1154 758 1158
rect 702 1143 704 1147
rect 716 1142 720 1154
rect 751 1150 755 1154
rect 745 1146 755 1150
rect 720 1138 725 1142
rect 778 1138 781 1142
rect 745 1106 870 1110
rect 745 1092 749 1106
rect 696 1085 698 1089
rect 739 1088 752 1092
rect 696 1077 698 1081
rect 710 1080 719 1084
rect 696 1069 698 1073
rect 710 1068 714 1080
rect 745 1076 749 1088
rect 739 1072 749 1076
rect 714 1064 719 1068
rect 782 1064 785 1068
rect 836 1033 848 1037
rect 745 1016 823 1020
rect 745 1010 749 1016
rect 819 1011 823 1016
rect 844 1019 848 1033
rect 866 1027 870 1106
rect 896 1035 900 1163
rect 1041 1118 1045 1500
rect 1190 1485 1194 1552
rect 1189 1484 1232 1485
rect 1193 1480 1232 1484
rect 1184 1471 1209 1476
rect 1149 1467 1188 1471
rect 1149 1403 1153 1467
rect 1192 1443 1196 1447
rect 1207 1443 1211 1447
rect 1192 1438 1211 1443
rect 1192 1434 1196 1438
rect 1160 1430 1164 1434
rect 1168 1403 1172 1410
rect 1184 1403 1188 1424
rect 1199 1419 1203 1438
rect 1207 1428 1211 1438
rect 1215 1441 1219 1447
rect 1227 1441 1232 1480
rect 1215 1437 1232 1441
rect 1303 1455 1309 1815
rect 1215 1428 1219 1437
rect 1212 1403 1216 1411
rect 1149 1399 1161 1403
rect 1168 1399 1216 1403
rect 1168 1396 1172 1399
rect 1160 1382 1164 1386
rect 1041 1114 1195 1118
rect 961 1069 1091 1073
rect 1191 1070 1195 1114
rect 961 1039 965 1069
rect 955 1035 968 1039
rect 896 1031 914 1035
rect 928 1027 941 1031
rect 866 1023 914 1027
rect 844 1015 914 1019
rect 928 1015 932 1027
rect 961 1023 965 1035
rect 955 1019 965 1023
rect 928 1011 941 1015
rect 696 1003 698 1007
rect 710 1006 719 1010
rect 745 1006 752 1010
rect 819 1007 914 1011
rect 696 995 698 999
rect 710 994 714 1006
rect 745 1002 749 1006
rect 739 998 749 1002
rect 880 999 914 1003
rect 928 999 932 1011
rect 961 1007 965 1019
rect 955 1003 965 1007
rect 696 987 698 991
rect 710 990 719 994
rect 696 979 698 983
rect 710 978 714 990
rect 745 986 749 998
rect 739 982 749 986
rect 714 974 719 978
rect 792 974 795 978
rect 880 942 884 999
rect 932 995 941 999
rect 1018 995 1021 999
rect 746 938 884 942
rect 746 923 750 938
rect 740 919 753 923
rect 697 915 699 919
rect 713 911 726 915
rect 697 907 699 911
rect 697 899 699 903
rect 713 899 717 911
rect 746 907 750 919
rect 740 903 750 907
rect 713 895 726 899
rect 697 891 699 895
rect 697 881 699 886
rect 713 883 717 895
rect 746 891 750 903
rect 740 887 750 891
rect 717 879 726 883
rect 803 879 806 883
rect 750 675 905 679
rect 750 663 754 675
rect 701 656 703 660
rect 715 659 724 663
rect 750 659 757 663
rect 701 648 703 652
rect 715 647 719 659
rect 750 655 754 659
rect 744 651 754 655
rect 719 643 724 647
rect 777 643 780 647
rect 744 605 875 609
rect 744 597 748 605
rect 695 590 697 594
rect 738 593 751 597
rect 695 582 697 586
rect 709 585 718 589
rect 695 574 697 578
rect 709 573 713 585
rect 744 581 748 593
rect 738 577 748 581
rect 713 569 718 573
rect 781 569 784 573
rect 744 515 748 521
rect 871 520 875 605
rect 901 528 905 675
rect 1087 617 1091 1069
rect 1189 1069 1232 1070
rect 1193 1065 1232 1069
rect 1184 1056 1209 1061
rect 1149 1052 1188 1056
rect 1149 988 1153 1052
rect 1192 1026 1196 1032
rect 1207 1026 1211 1032
rect 1192 1022 1211 1026
rect 1192 1019 1196 1022
rect 1160 1015 1164 1019
rect 1168 988 1172 995
rect 1184 988 1188 1009
rect 1199 999 1203 1022
rect 1207 1013 1211 1022
rect 1215 1026 1219 1032
rect 1227 1026 1232 1065
rect 1215 1022 1232 1026
rect 1303 1035 1309 1449
rect 1215 1013 1219 1022
rect 1212 988 1216 996
rect 1149 984 1161 988
rect 1168 984 1216 988
rect 1168 981 1172 984
rect 1160 967 1164 971
rect 1087 613 1199 617
rect 968 531 972 541
rect 901 524 921 528
rect 933 527 942 531
rect 968 527 975 531
rect 1195 530 1199 613
rect 1189 529 1232 530
rect 871 516 921 520
rect 933 515 937 527
rect 968 523 972 527
rect 1193 525 1232 529
rect 962 519 972 523
rect 695 508 697 512
rect 709 511 718 515
rect 744 511 751 515
rect 695 500 697 504
rect 709 499 713 511
rect 744 507 748 511
rect 853 508 921 512
rect 933 511 942 515
rect 738 503 748 507
rect 695 492 697 496
rect 709 495 718 499
rect 695 484 697 488
rect 709 483 713 495
rect 744 491 748 503
rect 895 500 921 504
rect 738 487 748 491
rect 713 479 718 483
rect 744 458 748 487
rect 791 479 794 483
rect 895 458 899 500
rect 933 499 937 511
rect 968 507 972 519
rect 1184 516 1209 521
rect 1149 512 1188 516
rect 962 503 972 507
rect 744 454 899 458
rect 907 492 921 496
rect 933 495 942 499
rect 745 428 749 437
rect 739 424 752 428
rect 696 420 698 424
rect 712 416 725 420
rect 696 412 698 416
rect 696 404 698 408
rect 712 404 716 416
rect 745 412 749 424
rect 739 408 749 412
rect 712 400 725 404
rect 696 396 698 400
rect 696 387 698 391
rect 712 388 716 400
rect 745 396 749 408
rect 739 392 749 396
rect 716 384 725 388
rect 745 367 749 392
rect 802 384 805 388
rect 907 367 911 492
rect 745 363 911 367
rect 917 336 921 488
rect 933 483 937 495
rect 968 491 972 503
rect 962 487 972 491
rect 937 479 942 483
rect 741 332 921 336
rect 741 324 745 332
rect 692 317 694 321
rect 706 320 715 324
rect 741 320 748 324
rect 692 309 694 313
rect 706 308 710 320
rect 741 316 745 320
rect 735 312 745 316
rect 692 301 694 305
rect 706 304 715 308
rect 692 293 694 297
rect 706 292 710 304
rect 741 300 745 312
rect 735 296 745 300
rect 706 288 715 292
rect 692 284 694 288
rect 692 275 694 279
rect 706 276 710 288
rect 741 284 745 296
rect 735 280 745 284
rect 710 272 715 276
rect 808 272 811 276
rect 968 140 972 487
rect 1035 479 1038 483
rect 1149 448 1153 512
rect 1192 486 1196 492
rect 1207 486 1211 492
rect 1192 482 1211 486
rect 1192 479 1196 482
rect 1160 475 1164 479
rect 1168 448 1172 455
rect 1184 448 1188 469
rect 1199 461 1203 482
rect 1207 473 1211 482
rect 1215 486 1219 492
rect 1227 486 1232 525
rect 1215 482 1232 486
rect 1215 473 1219 482
rect 1212 448 1216 456
rect 1149 444 1161 448
rect 1168 444 1216 448
rect 1303 459 1309 1030
rect 1168 441 1172 444
rect 1160 427 1164 431
rect 1303 169 1309 454
rect 1338 1841 1343 2099
rect 1472 2071 1475 2099
rect 1502 2071 1505 2099
rect 1513 2091 1524 2096
rect 1517 2083 1522 2091
rect 1521 2079 1522 2083
rect 1542 2071 1545 2099
rect 1568 2091 1572 2099
rect 1557 2075 1563 2078
rect 1560 2068 1563 2075
rect 1560 2064 1569 2068
rect 1491 2052 1495 2055
rect 1521 2051 1525 2055
rect 1564 2052 1569 2056
rect 1564 2051 1568 2052
rect 1521 2047 1568 2051
rect 1491 2042 1495 2047
rect 1521 2042 1525 2047
rect 1564 2045 1568 2047
rect 1584 2048 1588 2071
rect 1608 2075 1612 2099
rect 1616 2048 1620 2055
rect 1564 2041 1569 2045
rect 1584 2044 1609 2048
rect 1616 2044 1627 2048
rect 1584 2038 1588 2044
rect 1616 2041 1620 2044
rect 1475 2014 1479 2032
rect 1505 2014 1510 2032
rect 1568 2014 1572 2028
rect 1608 2014 1612 2031
rect 1469 2009 1622 2014
rect 1338 1837 1618 1841
rect 1622 1837 1626 1841
rect 1338 1474 1343 1837
rect 1472 1809 1475 1837
rect 1502 1809 1505 1837
rect 1513 1829 1524 1834
rect 1517 1821 1522 1829
rect 1521 1817 1522 1821
rect 1542 1809 1545 1837
rect 1568 1829 1572 1837
rect 1557 1813 1563 1816
rect 1560 1806 1563 1813
rect 1560 1802 1569 1806
rect 1491 1790 1495 1793
rect 1521 1789 1525 1793
rect 1564 1790 1569 1794
rect 1564 1789 1568 1790
rect 1521 1785 1568 1789
rect 1491 1780 1495 1785
rect 1521 1780 1525 1785
rect 1564 1783 1568 1785
rect 1584 1786 1588 1809
rect 1608 1813 1612 1837
rect 1616 1786 1620 1793
rect 1564 1779 1569 1783
rect 1584 1782 1609 1786
rect 1616 1782 1627 1786
rect 1584 1776 1588 1782
rect 1616 1779 1620 1782
rect 1475 1752 1479 1770
rect 1505 1752 1510 1770
rect 1568 1752 1572 1766
rect 1608 1752 1612 1769
rect 1467 1747 1622 1752
rect 1338 1470 1618 1474
rect 1622 1470 1626 1474
rect 1338 1056 1343 1470
rect 1472 1442 1475 1470
rect 1502 1442 1505 1470
rect 1513 1462 1524 1467
rect 1517 1454 1522 1462
rect 1521 1450 1522 1454
rect 1542 1442 1545 1470
rect 1568 1462 1572 1470
rect 1557 1446 1563 1449
rect 1560 1439 1563 1446
rect 1560 1435 1569 1439
rect 1491 1423 1495 1426
rect 1521 1422 1525 1426
rect 1564 1423 1569 1427
rect 1564 1422 1568 1423
rect 1521 1418 1568 1422
rect 1491 1413 1495 1418
rect 1521 1413 1525 1418
rect 1564 1416 1568 1418
rect 1584 1419 1588 1442
rect 1608 1446 1612 1470
rect 1616 1419 1620 1426
rect 1564 1412 1569 1416
rect 1584 1415 1609 1419
rect 1616 1415 1627 1419
rect 1584 1409 1588 1415
rect 1616 1412 1620 1415
rect 1475 1385 1479 1403
rect 1505 1385 1510 1403
rect 1568 1385 1572 1399
rect 1608 1385 1612 1402
rect 1467 1380 1475 1385
rect 1480 1380 1622 1385
rect 1338 1052 1618 1056
rect 1622 1052 1626 1056
rect 1338 480 1343 1052
rect 1472 1024 1475 1052
rect 1502 1024 1505 1052
rect 1513 1044 1524 1049
rect 1517 1036 1522 1044
rect 1521 1032 1522 1036
rect 1542 1024 1545 1052
rect 1568 1044 1572 1052
rect 1557 1028 1563 1031
rect 1560 1021 1563 1028
rect 1560 1017 1569 1021
rect 1491 1005 1495 1008
rect 1521 1004 1525 1008
rect 1564 1005 1569 1009
rect 1564 1004 1568 1005
rect 1521 1000 1568 1004
rect 1491 995 1495 1000
rect 1521 995 1525 1000
rect 1564 998 1568 1000
rect 1584 1001 1588 1024
rect 1608 1028 1612 1052
rect 1616 1001 1620 1008
rect 1564 994 1569 998
rect 1584 997 1609 1001
rect 1616 997 1627 1001
rect 1584 991 1588 997
rect 1616 994 1620 997
rect 1475 967 1479 985
rect 1505 967 1510 985
rect 1568 967 1572 981
rect 1608 967 1612 984
rect 1467 962 1474 967
rect 1480 962 1622 967
rect 1338 476 1618 480
rect 1622 476 1626 480
rect 1338 190 1343 476
rect 1472 448 1475 476
rect 1502 448 1505 476
rect 1513 468 1524 473
rect 1517 460 1522 468
rect 1521 456 1522 460
rect 1542 448 1545 476
rect 1568 468 1572 476
rect 1557 452 1563 455
rect 1560 445 1563 452
rect 1560 441 1569 445
rect 1491 429 1495 432
rect 1521 428 1525 432
rect 1564 429 1569 433
rect 1564 428 1568 429
rect 1521 424 1568 428
rect 1491 419 1495 424
rect 1521 419 1525 424
rect 1564 422 1568 424
rect 1584 425 1588 448
rect 1608 452 1612 476
rect 1616 425 1620 432
rect 1564 418 1569 422
rect 1584 421 1609 425
rect 1616 421 1627 425
rect 1584 415 1588 421
rect 1616 418 1620 421
rect 1475 391 1479 409
rect 1505 391 1510 409
rect 1568 391 1572 405
rect 1608 391 1612 408
rect 1467 386 1473 391
rect 1479 386 1622 391
rect 1338 186 1618 190
rect 1622 186 1626 190
rect 1472 158 1475 186
rect 1480 170 1484 173
rect 1502 158 1505 186
rect 1513 178 1524 183
rect 1517 170 1522 178
rect 1521 166 1522 170
rect 1542 158 1545 186
rect 1568 178 1572 186
rect 1557 162 1563 165
rect 1560 155 1563 162
rect 1560 151 1569 155
rect 968 137 1446 140
rect 1491 139 1495 142
rect 968 136 1475 137
rect 1442 133 1475 136
rect 1521 138 1525 142
rect 1564 139 1569 143
rect 1564 138 1568 139
rect 1521 134 1568 138
rect 1491 129 1495 134
rect 1521 129 1525 134
rect 1564 132 1568 134
rect 1584 135 1588 158
rect 1608 162 1612 186
rect 1616 135 1620 142
rect 1564 128 1569 132
rect 1584 131 1609 135
rect 1616 131 1627 135
rect 1584 125 1588 131
rect 1616 128 1620 131
rect 1475 101 1479 119
rect 1505 101 1510 119
rect 1568 101 1572 115
rect 1608 101 1612 118
rect 1467 96 1473 101
rect 1479 96 1622 101
rect 42 0 197 5
<< m2contact >>
rect 1303 2210 1309 2216
rect 261 2121 268 2128
rect 248 2088 253 2093
rect 317 2099 322 2104
rect 433 2157 438 2162
rect 384 2010 389 2015
rect 210 1976 215 1981
rect 264 1980 269 1985
rect 367 1969 372 1974
rect 398 1973 403 1978
rect 260 1835 267 1842
rect 251 1814 256 1819
rect 317 1816 322 1821
rect 440 2064 445 2069
rect 448 1973 453 1978
rect 456 1964 461 1969
rect 260 1697 267 1703
rect 217 1690 222 1695
rect 370 1681 375 1686
rect 405 1685 410 1690
rect 260 1513 267 1520
rect 249 1485 254 1490
rect 317 1487 322 1492
rect 263 1368 268 1373
rect 212 1343 219 1350
rect 374 1355 379 1360
rect 405 1359 410 1364
rect 260 1033 265 1038
rect 250 994 255 999
rect 315 998 320 1003
rect 215 871 220 876
rect 373 870 378 875
rect 404 874 409 879
rect 259 536 265 542
rect 238 504 243 509
rect 314 508 319 513
rect 259 389 264 394
rect 218 381 223 386
rect 373 384 378 389
rect 399 384 404 389
rect 202 34 207 39
rect 432 34 437 39
rect 464 1782 469 1787
rect 472 1685 477 1690
rect 480 1674 485 1679
rect 488 1453 493 1458
rect 496 1359 501 1364
rect 504 1349 509 1354
rect 512 997 517 1002
rect 520 874 525 879
rect 528 811 533 816
rect 536 473 541 478
rect 544 379 549 384
rect 552 320 557 325
rect 1191 2141 1196 2146
rect 709 2081 714 2087
rect 1162 2094 1167 2099
rect 1303 2082 1309 2089
rect 805 1984 810 1990
rect 706 1820 711 1826
rect 887 1795 892 1801
rect 706 1746 711 1752
rect 714 1546 719 1552
rect 1159 1798 1164 1803
rect 1332 1943 1338 1949
rect 1303 1815 1309 1822
rect 708 1472 713 1478
rect 896 1456 901 1462
rect 708 1382 713 1388
rect 716 1133 721 1138
rect 710 1059 715 1064
rect 1160 1438 1165 1443
rect 1303 1449 1309 1455
rect 710 969 715 974
rect 923 993 928 999
rect 713 873 718 879
rect 715 637 720 643
rect 709 563 714 569
rect 1159 1023 1164 1028
rect 1303 1030 1309 1035
rect 709 473 714 479
rect 712 378 717 384
rect 928 477 933 483
rect 706 266 711 272
rect 1159 483 1164 488
rect 1303 454 1309 459
rect 1303 164 1309 169
<< pm12contact >>
rect 67 2128 72 2133
rect 87 2128 92 2133
rect 159 2068 164 2073
rect 65 1990 70 1995
rect 85 1990 90 1995
rect 157 1930 162 1935
rect 65 1849 70 1854
rect 85 1849 90 1854
rect 157 1789 162 1794
rect 65 1707 70 1712
rect 85 1707 90 1712
rect 157 1647 162 1652
rect 65 1520 70 1525
rect 85 1520 90 1525
rect 157 1460 162 1465
rect 65 1378 70 1383
rect 85 1378 90 1383
rect 157 1318 162 1323
rect 65 1030 70 1035
rect 85 1030 90 1035
rect 157 970 162 975
rect 63 889 68 894
rect 83 889 88 894
rect 155 829 160 834
rect 63 540 68 545
rect 83 540 88 545
rect 155 480 160 485
rect 63 399 68 404
rect 83 399 88 404
rect 155 339 160 344
rect 63 70 68 75
rect 83 70 88 75
rect 155 10 160 15
rect 1488 2079 1493 2084
rect 1508 2079 1513 2084
rect 1580 2019 1585 2024
rect 1488 1817 1493 1822
rect 1508 1817 1513 1822
rect 1580 1757 1585 1762
rect 1488 1450 1493 1455
rect 1508 1450 1513 1455
rect 1580 1390 1585 1395
rect 1488 1032 1493 1037
rect 1508 1032 1513 1037
rect 1580 972 1585 977
rect 1488 456 1493 461
rect 1508 456 1513 461
rect 1580 396 1585 401
rect 1488 166 1493 171
rect 1508 166 1513 171
rect 1580 106 1585 111
<< metal2 >>
rect 14 2216 1309 2222
rect 14 2106 20 2216
rect 433 2171 1196 2176
rect 433 2162 438 2171
rect 1191 2146 1196 2171
rect 42 2138 70 2141
rect 42 2106 45 2138
rect 66 2135 70 2138
rect 66 2133 92 2135
rect 66 2132 67 2133
rect 72 2132 87 2133
rect 14 2100 45 2106
rect 219 2121 261 2126
rect 14 1980 20 2100
rect 42 2070 45 2100
rect 42 2068 159 2070
rect 42 2067 163 2068
rect 40 2000 68 2003
rect 40 1980 43 2000
rect 64 1997 68 2000
rect 64 1995 90 1997
rect 64 1994 65 1995
rect 70 1994 85 1995
rect 219 1986 224 2121
rect 14 1974 43 1980
rect 210 1981 224 1986
rect 248 1985 253 2088
rect 317 2068 321 2099
rect 850 2095 1162 2099
rect 653 2081 709 2086
rect 317 2064 440 2068
rect 653 2043 657 2081
rect 850 2043 854 2095
rect 1463 2089 1491 2092
rect 1463 2085 1466 2089
rect 1309 2082 1466 2085
rect 1487 2086 1491 2089
rect 1487 2084 1513 2086
rect 1487 2083 1488 2084
rect 653 2039 854 2043
rect 653 2015 657 2039
rect 1463 2021 1466 2082
rect 1493 2083 1508 2084
rect 1463 2019 1580 2021
rect 1463 2018 1584 2019
rect 389 2010 657 2015
rect 653 1989 657 2010
rect 653 1986 805 1989
rect 248 1980 264 1985
rect 14 1814 20 1974
rect 40 1932 43 1974
rect 403 1974 448 1978
rect 367 1947 372 1969
rect 400 1964 456 1969
rect 400 1947 405 1964
rect 367 1942 405 1947
rect 40 1930 157 1932
rect 40 1929 161 1930
rect 40 1859 68 1862
rect 40 1814 43 1859
rect 64 1856 68 1859
rect 64 1854 90 1856
rect 64 1853 65 1854
rect 70 1853 85 1854
rect 217 1837 260 1842
rect 14 1808 43 1814
rect 14 1685 20 1808
rect 40 1791 43 1808
rect 40 1789 157 1791
rect 40 1788 161 1789
rect 40 1717 68 1720
rect 40 1685 43 1717
rect 64 1714 68 1717
rect 64 1712 90 1714
rect 64 1711 65 1712
rect 70 1711 85 1712
rect 217 1695 222 1837
rect 653 1825 657 1986
rect 1115 1944 1332 1949
rect 653 1820 706 1825
rect 251 1797 255 1814
rect 247 1793 255 1797
rect 247 1701 251 1793
rect 317 1786 321 1816
rect 317 1782 464 1786
rect 653 1751 657 1820
rect 1115 1803 1120 1944
rect 1463 1827 1491 1830
rect 1463 1819 1466 1827
rect 1487 1824 1491 1827
rect 1487 1822 1513 1824
rect 1487 1821 1488 1822
rect 1309 1816 1466 1819
rect 1493 1821 1508 1822
rect 878 1796 887 1801
rect 878 1782 883 1796
rect 1112 1798 1159 1803
rect 1112 1782 1117 1798
rect 878 1777 1117 1782
rect 653 1746 706 1751
rect 247 1697 260 1701
rect 14 1679 43 1685
rect 410 1685 472 1690
rect 14 1493 20 1679
rect 40 1649 43 1679
rect 40 1647 157 1649
rect 40 1646 161 1647
rect 370 1634 375 1681
rect 653 1681 657 1746
rect 878 1681 883 1777
rect 1463 1759 1466 1816
rect 1463 1757 1580 1759
rect 1463 1756 1584 1757
rect 405 1674 480 1679
rect 653 1676 883 1681
rect 405 1634 410 1674
rect 370 1629 410 1634
rect 653 1549 657 1676
rect 653 1546 714 1549
rect 40 1530 68 1533
rect 40 1493 43 1530
rect 64 1527 68 1530
rect 64 1525 90 1527
rect 64 1524 65 1525
rect 70 1524 85 1525
rect 212 1513 260 1518
rect 14 1487 43 1493
rect 14 1359 20 1487
rect 40 1462 43 1487
rect 40 1460 157 1462
rect 40 1459 161 1460
rect 40 1388 68 1391
rect 40 1359 43 1388
rect 64 1385 68 1388
rect 64 1383 90 1385
rect 64 1382 65 1383
rect 70 1382 85 1383
rect 14 1353 43 1359
rect 14 1127 20 1353
rect 40 1320 43 1353
rect 212 1355 217 1513
rect 249 1481 254 1485
rect 249 1372 253 1481
rect 317 1458 322 1487
rect 653 1475 657 1546
rect 653 1472 708 1475
rect 317 1453 488 1458
rect 653 1385 657 1472
rect 887 1457 896 1462
rect 887 1419 891 1457
rect 1463 1460 1491 1463
rect 1463 1452 1466 1460
rect 1487 1457 1491 1460
rect 1487 1455 1513 1457
rect 1487 1454 1488 1455
rect 1309 1449 1466 1452
rect 1493 1454 1508 1455
rect 1123 1439 1160 1443
rect 1123 1419 1127 1439
rect 887 1415 1127 1419
rect 653 1382 708 1385
rect 249 1368 263 1372
rect 212 1350 219 1355
rect 410 1359 496 1364
rect 40 1318 157 1320
rect 40 1317 161 1318
rect 374 1302 379 1355
rect 403 1349 504 1354
rect 403 1302 408 1349
rect 374 1297 408 1302
rect 653 1302 657 1382
rect 887 1302 891 1415
rect 1463 1392 1466 1449
rect 1463 1390 1580 1392
rect 1463 1389 1584 1390
rect 653 1297 891 1302
rect 653 1136 657 1297
rect 653 1133 716 1136
rect 0 1122 20 1127
rect 14 1013 20 1122
rect 653 1062 657 1133
rect 653 1059 710 1062
rect 40 1040 68 1043
rect 40 1013 43 1040
rect 64 1037 68 1040
rect 64 1035 90 1037
rect 64 1034 65 1035
rect 70 1034 85 1035
rect 215 1033 260 1038
rect 14 1007 43 1013
rect 14 859 20 1007
rect 40 972 43 1007
rect 40 970 157 972
rect 40 969 161 970
rect 38 899 66 902
rect 38 859 41 899
rect 62 896 66 899
rect 62 894 88 896
rect 62 893 63 894
rect 68 893 83 894
rect 215 876 220 1033
rect 250 991 255 994
rect 251 882 254 991
rect 315 968 320 998
rect 343 997 512 1002
rect 343 968 348 997
rect 315 963 348 968
rect 653 972 657 1059
rect 1463 1042 1491 1045
rect 1463 1033 1466 1042
rect 1487 1039 1491 1042
rect 1487 1037 1513 1039
rect 1487 1036 1488 1037
rect 1309 1030 1466 1033
rect 1493 1036 1508 1037
rect 1119 1024 1159 1028
rect 911 994 923 998
rect 911 983 915 994
rect 1119 983 1123 1024
rect 911 979 1123 983
rect 653 969 710 972
rect 251 879 260 882
rect 409 874 520 879
rect 653 876 657 969
rect 14 853 42 859
rect 14 503 20 853
rect 38 831 41 853
rect 38 829 155 831
rect 38 828 159 829
rect 373 816 378 870
rect 653 873 713 876
rect 373 811 528 816
rect 653 798 657 873
rect 911 798 915 979
rect 1463 974 1466 1030
rect 1463 972 1580 974
rect 1463 971 1584 972
rect 653 794 915 798
rect 653 641 657 794
rect 653 637 715 641
rect 653 566 657 637
rect 653 563 709 566
rect 38 550 66 553
rect 38 503 41 550
rect 62 547 66 550
rect 62 545 88 547
rect 62 544 63 545
rect 68 544 83 545
rect 219 538 259 542
rect 14 497 42 503
rect 14 372 20 497
rect 38 482 41 497
rect 38 480 155 482
rect 38 479 159 480
rect 38 409 66 412
rect 38 372 41 409
rect 62 406 66 409
rect 62 404 88 406
rect 62 403 63 404
rect 68 403 83 404
rect 219 390 223 538
rect 218 386 223 390
rect 238 394 243 504
rect 314 478 319 508
rect 314 473 536 478
rect 653 476 657 563
rect 1110 483 1159 487
rect 653 473 709 476
rect 918 478 928 482
rect 238 389 259 394
rect 14 366 42 372
rect 14 49 20 366
rect 38 341 41 366
rect 38 339 155 341
rect 38 338 159 339
rect 373 325 378 384
rect 399 379 544 384
rect 653 381 657 473
rect 918 455 922 478
rect 1110 455 1114 483
rect 1463 466 1491 469
rect 918 451 1114 455
rect 1463 457 1466 466
rect 1487 463 1491 466
rect 1487 461 1513 463
rect 1487 460 1488 461
rect 1309 454 1466 457
rect 1493 460 1508 461
rect 653 378 712 381
rect 373 320 552 325
rect 653 269 657 378
rect 653 266 706 269
rect 653 182 657 266
rect 918 182 922 451
rect 1463 398 1466 454
rect 1463 396 1580 398
rect 1463 395 1584 396
rect 653 178 922 182
rect 1463 176 1491 179
rect 1463 167 1466 176
rect 1487 173 1491 176
rect 1487 171 1513 173
rect 1487 170 1488 171
rect 1309 164 1466 167
rect 1493 170 1508 171
rect 1463 108 1466 164
rect 1463 106 1580 108
rect 1463 105 1584 106
rect 38 80 66 83
rect 38 49 41 80
rect 62 77 66 80
rect 62 75 88 77
rect 62 74 63 75
rect 68 74 83 75
rect 14 43 42 49
rect 38 12 41 43
rect 207 34 432 39
rect 38 10 155 12
rect 38 9 159 10
<< m3contact >>
rect 125 547 130 552
<< m123contact >>
rect 204 2148 209 2153
rect 87 2140 92 2145
rect 129 2138 134 2143
rect 1145 2122 1151 2129
rect 70 2096 75 2101
rect 202 2010 207 2015
rect 85 2002 90 2007
rect 127 1997 132 2002
rect 274 2112 279 2117
rect 441 2101 446 2106
rect 691 2101 696 2106
rect 433 2090 438 2095
rect 691 2090 696 2095
rect 771 2082 776 2087
rect 565 2069 570 2074
rect 1508 2091 1513 2096
rect 1550 2086 1555 2091
rect 1200 2067 1205 2072
rect 1161 2034 1166 2039
rect 1471 2045 1476 2050
rect 1491 2047 1496 2052
rect 375 2008 380 2013
rect 457 1994 462 1999
rect 1463 2007 1469 2014
rect 786 1994 791 1999
rect 565 1980 570 1985
rect 276 1966 281 1971
rect 68 1958 73 1963
rect 202 1869 207 1874
rect 85 1861 90 1866
rect 127 1856 132 1861
rect 68 1817 73 1822
rect 202 1727 207 1732
rect 85 1719 90 1724
rect 127 1714 132 1719
rect 465 1840 470 1845
rect 274 1829 279 1834
rect 449 1829 454 1834
rect 867 1985 872 1990
rect 687 1840 692 1845
rect 687 1829 692 1834
rect 768 1821 773 1826
rect 565 1811 570 1816
rect 481 1795 486 1801
rect 465 1773 470 1778
rect 441 1765 446 1770
rect 433 1756 438 1761
rect 858 1810 864 1816
rect 1142 1823 1149 1828
rect 1508 1829 1513 1834
rect 1550 1824 1555 1829
rect 964 1792 969 1797
rect 681 1774 686 1779
rect 681 1765 686 1770
rect 681 1756 686 1761
rect 772 1747 777 1752
rect 565 1737 570 1742
rect 378 1721 383 1726
rect 276 1683 281 1688
rect 68 1675 73 1680
rect 1198 1772 1203 1777
rect 1470 1784 1475 1789
rect 1491 1785 1496 1790
rect 1461 1747 1467 1752
rect 1159 1733 1164 1738
rect 489 1564 494 1569
rect 473 1554 478 1559
rect 695 1565 700 1570
rect 695 1555 700 1560
rect 776 1547 781 1552
rect 202 1540 207 1545
rect 85 1532 90 1537
rect 565 1533 570 1538
rect 127 1527 132 1532
rect 68 1488 73 1493
rect 202 1398 207 1403
rect 85 1390 90 1395
rect 127 1385 132 1390
rect 274 1500 279 1505
rect 489 1499 494 1504
rect 465 1490 470 1495
rect 449 1481 454 1486
rect 689 1500 694 1505
rect 689 1491 694 1496
rect 689 1482 694 1487
rect 780 1473 785 1478
rect 565 1463 570 1468
rect 505 1449 510 1454
rect 489 1417 494 1422
rect 465 1408 470 1413
rect 441 1399 446 1404
rect 378 1394 383 1399
rect 433 1390 438 1395
rect 1142 1464 1149 1469
rect 848 1448 854 1454
rect 689 1418 694 1423
rect 1508 1462 1513 1467
rect 983 1453 988 1458
rect 1550 1457 1555 1462
rect 689 1409 694 1414
rect 689 1400 694 1405
rect 689 1391 694 1396
rect 790 1383 795 1388
rect 565 1373 570 1378
rect 68 1346 73 1351
rect 276 1354 281 1359
rect 1198 1414 1203 1419
rect 1470 1417 1475 1422
rect 1491 1418 1496 1423
rect 1475 1380 1480 1385
rect 1159 1373 1164 1378
rect 513 1151 518 1156
rect 497 1142 502 1147
rect 697 1152 702 1157
rect 697 1143 702 1148
rect 778 1133 783 1138
rect 565 1128 570 1133
rect 513 1085 518 1090
rect 489 1076 494 1081
rect 473 1067 478 1073
rect 691 1086 696 1091
rect 691 1077 696 1082
rect 691 1068 696 1073
rect 782 1059 787 1064
rect 202 1050 207 1055
rect 565 1049 570 1054
rect 85 1042 90 1047
rect 127 1037 132 1042
rect 68 998 73 1003
rect 200 909 205 914
rect 83 901 88 906
rect 125 896 130 901
rect 529 1032 534 1038
rect 513 1020 518 1026
rect 274 1011 279 1016
rect 489 1008 494 1013
rect 465 985 470 991
rect 449 976 454 981
rect 1142 1047 1149 1052
rect 1508 1044 1513 1049
rect 831 1032 836 1038
rect 1550 1039 1555 1044
rect 691 1004 696 1009
rect 691 995 696 1000
rect 691 986 696 991
rect 1018 990 1023 995
rect 1198 994 1203 999
rect 691 977 696 982
rect 792 969 797 974
rect 565 959 570 964
rect 513 915 518 920
rect 377 909 382 914
rect 489 906 494 911
rect 432 900 437 906
rect 465 897 470 902
rect 441 888 446 893
rect 692 916 697 921
rect 692 907 697 912
rect 692 898 697 903
rect 692 889 697 894
rect 692 880 697 885
rect 274 865 279 870
rect 66 857 71 862
rect 803 874 808 879
rect 565 864 570 869
rect 1470 999 1475 1004
rect 1491 1000 1496 1005
rect 1159 958 1164 963
rect 1474 962 1480 967
rect 537 655 542 660
rect 521 646 526 651
rect 696 656 701 661
rect 696 647 701 652
rect 777 638 782 643
rect 565 628 570 633
rect 537 590 542 595
rect 513 581 518 586
rect 497 572 502 577
rect 690 591 695 596
rect 690 582 695 587
rect 690 573 695 578
rect 200 560 205 565
rect 781 564 786 569
rect 83 552 88 557
rect 565 554 570 559
rect 66 508 71 513
rect 200 419 205 424
rect 83 411 88 416
rect 125 406 130 411
rect 553 538 558 543
rect 274 521 279 526
rect 537 508 542 513
rect 513 499 518 504
rect 489 490 494 495
rect 472 485 478 490
rect 690 509 695 514
rect 848 508 853 513
rect 690 500 695 505
rect 1142 504 1149 509
rect 690 491 695 496
rect 690 482 695 487
rect 791 474 796 479
rect 565 464 570 469
rect 377 423 382 428
rect 537 420 542 425
rect 513 411 518 416
rect 489 402 494 407
rect 449 394 454 400
rect 465 393 470 398
rect 273 375 278 380
rect 66 367 71 372
rect 1035 474 1040 479
rect 1508 468 1513 473
rect 1198 456 1203 461
rect 1550 463 1555 468
rect 691 421 696 426
rect 691 412 696 417
rect 691 403 696 408
rect 691 394 696 399
rect 691 385 696 390
rect 802 379 807 384
rect 565 369 570 374
rect 537 311 542 316
rect 513 302 518 307
rect 489 293 494 298
rect 441 283 446 288
rect 465 284 470 289
rect 433 267 438 272
rect 687 318 692 323
rect 687 309 692 314
rect 687 300 692 305
rect 687 291 692 296
rect 687 282 692 287
rect 687 273 692 278
rect 808 267 813 272
rect 565 257 570 262
rect 1159 418 1164 423
rect 1470 423 1475 428
rect 1491 424 1496 429
rect 1473 386 1479 391
rect 1508 178 1513 183
rect 1550 173 1555 178
rect 1491 134 1496 139
rect 1473 96 1479 101
rect 200 90 205 95
rect 83 82 88 87
rect 125 77 130 82
rect 66 38 71 43
<< metal3 >>
rect 117 2200 1534 2203
rect 77 2140 87 2145
rect 117 2141 120 2200
rect 209 2148 232 2152
rect 77 2101 80 2140
rect 117 2138 129 2141
rect 75 2096 81 2101
rect 75 2002 85 2007
rect 75 1963 78 2002
rect 117 2000 120 2138
rect 228 2117 232 2148
rect 691 2124 1145 2129
rect 228 2112 274 2117
rect 228 2014 232 2112
rect 691 2106 696 2124
rect 446 2101 691 2104
rect 438 2090 691 2093
rect 1498 2091 1508 2096
rect 771 2073 775 2082
rect 570 2069 775 2073
rect 1200 2048 1205 2067
rect 1498 2052 1501 2091
rect 1531 2090 1534 2200
rect 1531 2087 1550 2090
rect 1200 2043 1471 2048
rect 1496 2047 1502 2052
rect 207 2013 232 2014
rect 207 2010 375 2013
rect 228 2009 375 2010
rect 117 1997 127 2000
rect 73 1958 79 1963
rect 75 1861 85 1866
rect 75 1822 78 1861
rect 117 1859 120 1997
rect 228 1971 232 2009
rect 462 1994 786 1997
rect 1161 1985 1166 2034
rect 1269 2010 1463 2015
rect 1269 1985 1274 2010
rect 570 1980 1274 1985
rect 228 1966 276 1971
rect 228 1873 232 1966
rect 207 1869 232 1873
rect 117 1856 127 1859
rect 73 1817 79 1822
rect 75 1719 85 1724
rect 75 1680 78 1719
rect 117 1717 120 1856
rect 228 1834 232 1869
rect 670 1869 1021 1872
rect 670 1843 673 1869
rect 470 1840 687 1843
rect 228 1829 274 1834
rect 454 1829 687 1832
rect 228 1731 232 1829
rect 1018 1828 1021 1869
rect 1498 1829 1508 1834
rect 1018 1825 1142 1828
rect 768 1816 773 1821
rect 570 1811 773 1816
rect 834 1810 858 1816
rect 834 1801 840 1810
rect 486 1795 840 1801
rect 470 1774 681 1777
rect 446 1765 681 1768
rect 438 1756 681 1759
rect 772 1742 777 1747
rect 964 1742 969 1792
rect 1498 1790 1501 1829
rect 1531 1828 1534 2087
rect 1531 1825 1550 1828
rect 1255 1784 1470 1789
rect 1496 1785 1502 1790
rect 1198 1757 1203 1772
rect 1255 1757 1260 1784
rect 1198 1752 1260 1757
rect 1455 1747 1461 1752
rect 570 1738 1118 1742
rect 570 1737 1159 1738
rect 1113 1733 1159 1737
rect 207 1727 232 1731
rect 228 1726 232 1727
rect 228 1722 378 1726
rect 117 1714 127 1717
rect 73 1675 79 1680
rect 75 1532 85 1537
rect 75 1493 78 1532
rect 117 1530 120 1714
rect 228 1688 232 1722
rect 1150 1720 1155 1733
rect 1455 1720 1460 1747
rect 1150 1715 1460 1720
rect 228 1683 276 1688
rect 228 1544 232 1683
rect 686 1623 913 1626
rect 686 1568 689 1623
rect 494 1565 695 1568
rect 910 1560 913 1623
rect 478 1555 695 1558
rect 910 1557 975 1560
rect 207 1540 232 1544
rect 117 1527 127 1530
rect 73 1488 79 1493
rect 75 1390 85 1395
rect 75 1351 78 1390
rect 117 1388 120 1527
rect 228 1505 232 1540
rect 776 1538 781 1547
rect 570 1533 781 1538
rect 972 1525 975 1557
rect 972 1522 1086 1525
rect 228 1500 274 1505
rect 228 1402 232 1500
rect 494 1500 689 1503
rect 470 1491 689 1494
rect 454 1482 689 1485
rect 780 1468 785 1473
rect 570 1463 785 1468
rect 1083 1467 1086 1522
rect 1083 1464 1142 1467
rect 1498 1462 1508 1467
rect 510 1449 848 1453
rect 494 1418 689 1421
rect 470 1409 689 1412
rect 207 1399 232 1402
rect 446 1400 689 1403
rect 207 1398 378 1399
rect 228 1395 378 1398
rect 117 1385 127 1388
rect 73 1346 79 1351
rect 117 1177 120 1385
rect 228 1359 232 1395
rect 438 1391 689 1394
rect 790 1380 795 1383
rect 983 1380 988 1453
rect 1498 1423 1501 1462
rect 1531 1461 1534 1825
rect 1531 1458 1550 1461
rect 1198 1389 1203 1414
rect 1440 1417 1470 1422
rect 1496 1418 1502 1423
rect 1440 1389 1445 1417
rect 1198 1384 1445 1389
rect 790 1378 1096 1380
rect 570 1377 1096 1378
rect 570 1375 1159 1377
rect 570 1373 795 1375
rect 1091 1372 1159 1375
rect 228 1354 276 1359
rect 1138 1357 1143 1372
rect 1475 1357 1480 1380
rect 228 1218 232 1354
rect 1138 1352 1480 1357
rect 223 1214 232 1218
rect 105 1173 120 1177
rect 75 1042 85 1047
rect 75 1003 78 1042
rect 117 1040 120 1173
rect 228 1054 232 1214
rect 688 1195 1016 1198
rect 688 1155 691 1195
rect 518 1152 697 1155
rect 502 1143 697 1146
rect 570 1128 783 1133
rect 518 1086 691 1089
rect 494 1077 691 1080
rect 478 1068 691 1071
rect 782 1054 787 1059
rect 207 1050 232 1054
rect 117 1037 127 1040
rect 73 998 79 1003
rect 73 901 83 906
rect 73 862 76 901
rect 117 899 120 1037
rect 228 1016 232 1050
rect 570 1049 787 1054
rect 1013 1052 1016 1195
rect 1013 1049 1142 1052
rect 1498 1044 1508 1049
rect 534 1032 831 1038
rect 518 1021 571 1024
rect 228 1011 274 1016
rect 228 914 232 1011
rect 494 1009 560 1012
rect 557 998 560 1009
rect 568 1007 571 1021
rect 568 1004 691 1007
rect 1498 1005 1501 1044
rect 1531 1043 1534 1458
rect 1531 1040 1550 1043
rect 557 995 691 998
rect 470 986 691 989
rect 454 977 691 980
rect 792 968 797 969
rect 1018 968 1023 990
rect 1198 977 1203 994
rect 1444 997 1470 1002
rect 1496 1000 1502 1005
rect 1444 977 1449 997
rect 1198 972 1449 977
rect 792 964 1124 968
rect 570 963 1124 964
rect 570 959 797 963
rect 1119 958 1159 963
rect 1148 926 1153 958
rect 1474 926 1479 962
rect 1148 921 1479 926
rect 518 916 692 919
rect 228 913 377 914
rect 205 910 377 913
rect 205 909 232 910
rect 117 896 125 899
rect 71 857 77 862
rect 73 552 83 557
rect 73 513 76 552
rect 117 550 120 896
rect 228 870 232 909
rect 494 907 692 910
rect 434 883 437 900
rect 470 898 692 901
rect 446 889 692 892
rect 434 880 692 883
rect 228 865 274 870
rect 803 869 808 874
rect 228 564 232 865
rect 570 864 808 869
rect 682 717 1005 720
rect 682 659 685 717
rect 542 656 696 659
rect 526 647 696 650
rect 777 633 782 638
rect 570 628 786 633
rect 542 591 690 594
rect 518 582 690 585
rect 1002 585 1005 717
rect 1002 582 1102 585
rect 502 573 690 576
rect 205 560 232 564
rect 117 547 125 550
rect 71 508 77 513
rect 73 411 83 416
rect 73 372 76 411
rect 117 409 120 547
rect 228 526 232 560
rect 781 559 786 564
rect 570 554 794 559
rect 558 538 848 543
rect 228 521 274 526
rect 228 428 232 521
rect 542 509 690 512
rect 843 508 848 538
rect 1099 508 1102 582
rect 1099 505 1142 508
rect 518 500 690 503
rect 494 491 690 494
rect 473 482 690 485
rect 791 469 796 474
rect 1035 469 1040 474
rect 570 464 1040 469
rect 1498 468 1508 473
rect 228 424 377 428
rect 228 423 232 424
rect 205 419 232 423
rect 542 421 691 424
rect 1033 422 1038 464
rect 1198 427 1203 456
rect 1498 429 1501 468
rect 1531 467 1534 1040
rect 1531 464 1550 467
rect 117 406 125 409
rect 71 367 77 372
rect 73 82 83 87
rect 73 43 76 82
rect 117 80 120 406
rect 228 380 232 419
rect 1033 417 1159 422
rect 1198 422 1470 427
rect 1496 424 1502 429
rect 518 412 691 415
rect 494 403 691 406
rect 449 388 452 394
rect 470 394 691 397
rect 449 385 691 388
rect 228 375 273 380
rect 228 94 232 375
rect 802 374 807 379
rect 1149 383 1154 417
rect 1473 383 1478 386
rect 1149 378 1478 383
rect 570 369 807 374
rect 569 318 687 321
rect 569 315 572 318
rect 542 312 572 315
rect 576 309 687 312
rect 576 306 579 309
rect 518 303 579 306
rect 583 300 687 303
rect 583 297 586 300
rect 494 294 586 297
rect 591 291 687 294
rect 591 288 594 291
rect 470 285 594 288
rect 441 279 444 283
rect 598 282 687 285
rect 598 279 601 282
rect 441 276 601 279
rect 607 273 687 276
rect 607 271 610 273
rect 438 268 610 271
rect 808 262 813 267
rect 570 257 813 262
rect 205 90 232 94
rect 1247 93 1252 378
rect 1498 178 1508 183
rect 1498 139 1501 178
rect 1531 177 1534 464
rect 1531 174 1550 177
rect 1496 134 1502 139
rect 1473 93 1478 96
rect 1247 88 1478 93
rect 1531 85 1534 174
rect 117 77 125 80
rect 71 38 77 43
<< metal4 >>
rect 479 2087 483 2091
<< labels >>
rlabel metal1 59 2132 63 2135 1 a0
rlabel metal1 57 1994 61 1997 1 b0
rlabel metal1 57 1853 61 1856 1 a1
rlabel metal1 57 1711 61 1714 1 b1
rlabel metal1 57 1524 61 1527 1 a2
rlabel metal1 57 1382 61 1385 1 b2
rlabel metal1 57 1034 61 1037 1 a3
rlabel metal1 55 893 59 896 1 b3
rlabel metal1 55 544 59 547 1 a4
rlabel metal1 55 403 59 406 1 b4
rlabel metal1 55 74 59 77 1 c0
rlabel metal2 0 1122 14 1127 1 clk
rlabel metal3 105 1173 117 1177 1 rst
rlabel metal1 33 676 38 680 1 gnd
rlabel metal3 223 1214 228 1218 1 vdd
rlabel metal1 177 2093 180 2097 1 qb0
rlabel metal1 201 2093 204 2097 1 q0
rlabel metal1 178 1955 181 1959 1 qb5
rlabel metal1 200 1955 203 1959 1 q5
rlabel metal1 180 1814 183 1818 1 qb1
rlabel metal1 200 1814 203 1818 1 q1
rlabel metal1 175 1672 178 1676 1 qb6
rlabel metal1 200 1672 203 1676 1 q6
rlabel metal1 176 1485 179 1489 1 qb2
rlabel metal1 199 1485 202 1489 1 q2
rlabel metal1 176 1343 179 1347 1 qb7
rlabel metal1 199 1343 202 1347 1 q7
rlabel metal1 177 995 180 999 1 qb3
rlabel metal1 199 995 202 999 1 q3
rlabel metal1 175 854 178 858 1 qb8
rlabel metal1 197 854 200 858 1 q8
rlabel metal1 177 505 180 509 1 qb4
rlabel metal1 197 505 200 509 1 q4
rlabel metal1 176 364 179 368 1 qb9
rlabel metal1 197 364 200 368 1 q9
rlabel metal1 197 35 200 39 1 qc0
rlabel metal1 174 35 177 39 1 qbc0
rlabel metal1 317 2104 321 2108 1 p0
rlabel metal1 367 1974 370 1978 1 g0_bar
rlabel metal1 395 1974 398 1978 1 g0
rlabel metal1 317 1821 320 1825 1 p1
rlabel metal1 371 1686 374 1690 1 g1_bar
rlabel metal1 401 1686 404 1690 1 g1
rlabel metal1 317 1492 320 1496 1 p2
rlabel metal1 377 1360 380 1364 1 g2_bar
rlabel metal1 397 1360 400 1364 1 g2
rlabel metal1 315 1003 318 1007 1 p3
rlabel metal1 376 875 379 879 1 g3_bar
rlabel metal1 398 875 401 879 1 g3
rlabel metal1 314 513 317 517 1 p4
rlabel metal1 376 389 379 393 1 g4_bar
rlabel metal1 401 389 404 393 1 g4
rlabel metal1 840 2016 844 2019 1 c1
rlabel metal1 927 1831 931 1834 1 c2
rlabel metal1 936 1501 940 1504 1 c3
rlabel metal1 961 1046 965 1048 1 c4
rlabel metal1 968 539 972 541 1 cout
rlabel metal1 1201 2086 1205 2089 1 s0
rlabel metal1 1199 1790 1203 1793 1 s1
rlabel metal1 1199 1015 1203 1018 1 s3
rlabel metal1 1199 475 1203 478 1 s4
rlabel metal1 1600 2044 1604 2048 1 qbs0
rlabel metal1 1623 2044 1627 2048 7 qs0
rlabel metal1 1601 1782 1605 1786 1 qbs1
rlabel metal1 1623 1782 1627 1786 7 qs1
rlabel metal1 1623 1415 1627 1419 7 qs2
rlabel metal1 1602 1415 1606 1419 1 qbs2
rlabel metal1 1604 997 1608 1001 1 qbs3
rlabel metal1 1622 997 1626 1001 7 qs3
rlabel metal1 1623 421 1627 425 7 qs4
rlabel metal1 1199 1433 1203 1438 1 s2
rlabel metal1 1623 131 1626 135 7 qcout
rlabel metal1 1600 131 1603 135 1 qbcout
rlabel metal1 1603 421 1607 425 1 qbs4
<< end >>
