magic
tech scmos
timestamp 1763396525
<< nwell >>
rect 9 -76 49 -12
<< ntransistor >>
rect 56 -25 116 -23
rect 56 -33 116 -31
rect 56 -41 116 -39
rect 56 -49 116 -47
rect 56 -57 116 -55
rect 56 -65 116 -63
<< ptransistor >>
rect 23 -25 43 -23
rect 23 -33 43 -31
rect 23 -41 43 -39
rect 23 -49 43 -47
rect 23 -57 43 -55
rect 23 -65 43 -63
<< ndiffusion >>
rect 56 -23 116 -22
rect 56 -26 116 -25
rect 56 -31 116 -30
rect 56 -34 116 -33
rect 56 -39 116 -38
rect 56 -42 116 -41
rect 56 -47 116 -46
rect 56 -50 116 -49
rect 56 -55 116 -54
rect 56 -58 116 -57
rect 56 -63 116 -62
rect 56 -66 116 -65
<< pdiffusion >>
rect 23 -23 43 -22
rect 23 -26 43 -25
rect 23 -31 43 -30
rect 23 -34 43 -33
rect 23 -39 43 -38
rect 23 -42 43 -41
rect 23 -47 43 -46
rect 23 -50 43 -49
rect 23 -55 43 -54
rect 23 -58 43 -57
rect 23 -63 43 -62
rect 23 -66 43 -65
<< ndcontact >>
rect 56 -22 116 -18
rect 56 -30 116 -26
rect 56 -38 116 -34
rect 56 -46 116 -42
rect 56 -54 116 -50
rect 56 -62 116 -58
rect 56 -70 116 -66
<< pdcontact >>
rect 23 -22 43 -18
rect 23 -30 43 -26
rect 23 -38 43 -34
rect 23 -46 43 -42
rect 23 -54 43 -50
rect 23 -62 43 -58
rect 23 -70 43 -66
<< psubstratepcontact >>
rect 121 -70 125 -66
<< nsubstratencontact >>
rect 14 -70 18 -66
<< polysilicon >>
rect 6 -25 23 -23
rect 43 -25 56 -23
rect 116 -25 119 -23
rect 6 -33 23 -31
rect 43 -33 56 -31
rect 116 -33 119 -31
rect 6 -41 23 -39
rect 43 -41 56 -39
rect 116 -41 119 -39
rect 6 -49 23 -47
rect 43 -49 56 -47
rect 116 -49 119 -47
rect 6 -57 23 -55
rect 43 -57 56 -55
rect 116 -57 119 -55
rect 6 -65 23 -63
rect 43 -65 56 -63
rect 116 -65 119 -63
<< polycontact >>
rect 2 -25 6 -21
rect 2 -33 6 -29
rect 2 -41 6 -37
rect 2 -49 6 -45
rect 2 -57 6 -53
rect 2 -65 6 -61
<< metal1 >>
rect 49 -18 53 -8
rect 0 -25 2 -21
rect 14 -22 23 -18
rect 49 -22 56 -18
rect 0 -33 2 -29
rect 14 -34 18 -22
rect 49 -26 53 -22
rect 43 -30 53 -26
rect 0 -41 2 -37
rect 14 -38 23 -34
rect 0 -49 2 -45
rect 14 -50 18 -38
rect 49 -42 53 -30
rect 43 -46 53 -42
rect 0 -57 2 -53
rect 14 -54 23 -50
rect 0 -65 2 -61
rect 14 -66 18 -54
rect 49 -58 53 -46
rect 43 -62 53 -58
rect 18 -70 23 -66
rect 116 -70 121 -66
<< labels >>
rlabel metal1 0 -65 2 -63 3 a
rlabel metal1 0 -57 2 -55 3 b
rlabel metal1 0 -49 2 -47 3 c
rlabel metal1 0 -41 2 -39 3 d
rlabel metal1 0 -33 2 -31 3 e
rlabel metal1 0 -25 2 -23 3 f
rlabel psubstratepcontact 121 -70 125 -66 7 gnd
rlabel nsubstratencontact 14 -70 18 -66 7 vdd
rlabel metal1 49 -11 53 -8 5 vo
<< end >>
