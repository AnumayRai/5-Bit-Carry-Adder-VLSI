D Flip Flop
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

.param width_P= {20*lambda}
.param width_N= {10*lambda}
    
Vdd	vdd	gnd	'SUPPLY'
vclk clk gnd pulse 0 1.8 0ns 0ns 0ns 5ns 10ns
vin d gnd pulse 0 1.8 2ns 0ns 0ns 20ns 40ns
vrst rst gnd pulse 1.8 0 80ns 0ns 0ns 5ns 100ns
.option scale=0.09u

M1000 a clk a_13_6# vdd cmosp w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1001 a d gnd Gnd cmosn w=10 l=2
+  ad=130 pd=46 as=200 ps=120
M1002 qb b vdd vdd cmosp w=20 l=2
+  ad=260 pd=66 as=500 ps=250
M1003 q qb vdd vdd cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1004 b a a_43_n17# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=60 ps=32
M1005 a_43_n17# clk gnd Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 q qb gnd Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1007 a_13_6# d vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_106_n21# b gnd Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1009 qb clk a_106_n21# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1010 b a a_43_6# vdd cmosp w=20 l=2
+  ad=200 pd=100 as=120 ps=52
M1011 b rst vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 a_43_6# clk vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd q 0.25fF
C1 rst vdd 0.15fF
C2 gnd b 0.05fF
C3 a_43_n17# b 0.10fF
C4 vdd d 0.19fF
C5 d clk 0.10fF
C6 vdd clk 1.04fF
C7 rst b 0.01fF
C8 a_43_6# vdd 0.21fF
C9 gnd qb 0.05fF
C10 a_13_6# a 0.21fF
C11 qb q 0.05fF
C12 gnd a_106_n21# 0.10fF
C13 vdd b 0.80fF
C14 b clk 0.03fF
C15 a_43_6# b 0.21fF
C16 qb vdd 0.41fF
C17 qb clk 0.01fF
C18 gnd a 0.10fF
C19 a_13_6# d 0.01fF
C20 vdd a_13_6# 0.21fF
C21 vdd a 0.77fF
C22 a clk 0.27fF
C23 gnd a_43_n17# 0.10fF
C24 gnd q 0.10fF
C25 qb a_106_n21# 0.10fF
C26 a b 0.01fF
C27 gnd clk 0.32fF
C28 a_106_n21# Gnd 0.01fF
C29 a_43_n17# Gnd 0.01fF
C30 gnd Gnd 0.47fF
C31 q Gnd 0.06fF
C32 qb Gnd 0.23fF
C33 a Gnd 0.09fF
C34 clk Gnd 0.10fF
C35 d Gnd 0.08fF
C36 b Gnd 0.08fF
C37 vdd Gnd 3.43fF

.tran 0.1n 200n

.measure tran tcq
+TRIG v(d) VAL=0.9 RISE=1
+TARG v(q) VAL=0.9 RISE=1

.measure tran SetupTime
+TRIG v(d) VAL=0.9 RISE=1
+TARG v(a) VAL=0.9 FALL=1

.measure tran HoldTime
+TRIG v(a) VAL=0.9 RISE=1
+TARG v(b) VAL=0.9 FALL=1

.control
set hcopypscolor = 1 *White background for saving plots
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7))
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7))


run
plot v(clk)+8  v(rst)+6 v(d)+4 v(q)+2 

.endc
.end
