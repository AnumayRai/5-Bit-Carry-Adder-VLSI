2 input XOR
.include TSMC_180nm.txt

.param SUPPLY = 1.8
.param LAMBDA = 0.09u
.param width_P= {20*lambda}
.param width_N= {10*lambda}

.global gnd vdd

Vdd vdd gnd {SUPPLY}
Vin1  a   gnd PULSE(0 {SUPPLY} 0n 0n 0n 20n 40n)
Vin2  b   gnd PULSE(0 {SUPPLY} 0n 0n 0n 40n 80n)


Ma1 a_bar a vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

Ma2 a_bar a gnd gnd CMOSN W={width_N} L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M1 vo b a vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M2 vo b a_bar gnd CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

M3 vo a b vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

M4 vo a_bar b gnd CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}

.tran 0.1n 200n

.control
set hcopypscolor=1
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=green
set color5=orange
run
plot v(a)+8 v(b)+6 v(a_bar)+4  v(vo)
.endc
.end

