3-I/P NAND GATE
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

.param width_P= {20*lambda}
.param width_N= {3*10*lambda}
    
Vdd	vdd	gnd	'SUPPLY'
va a gnd pulse 0 1.8 2ns 0ns 0ns 20ns 40ns
vb b gnd pulse 0 1.8 1ns 0ns 0ns 40ns 80ns
vc c gnd pulse 0 1.8 0ns 0ns 0ns 80ns 160ns
.option scale=0.09u

M1000 vo a vdd vdd cmosp w=20 l=2
+  ad=220 pd=102 as=220 ps=102
M1001 vo c a_56_n25# Gnd cmosn w=30 l=2
+  ad=150 pd=70 as=180 ps=72
M1002 a_56_n25# b a_56_n33# Gnd cmosn w=30 l=2
+  ad=0 pd=0 as=180 ps=72
M1003 vo c vdd vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_56_n33# a gnd Gnd cmosn w=30 l=2
+  ad=0 pd=0 as=150 ps=70
M1005 vdd b vo vdd cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vo b 0.08fF
C1 a b 0.21fF
C2 vdd c 0.12fF
C3 c vo 0.08fF
C4 vdd vo 0.76fF
C5 gnd a_56_n33# 0.31fF
C6 a_56_n25# vo 0.36fF
C7 c b 0.21fF
C8 a_56_n25# a_56_n33# 0.31fF
C9 vdd b 0.20fF
C10 vo a_56_n33# 0.05fF
C11 a vdd 0.20fF

.tran 0.1n 200n

.control
set hcopypscolor = 1
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=green
set color5=orange
run
plot v(a)+6 v(b)+4 v(c)+2 v(vo)
.endc

.end
